interface aes_interface_inner;




endinterface
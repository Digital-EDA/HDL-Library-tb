
module rot (
        input         clka,
        input         rsta,
        input  [8:0]  addra,
        output [31:0] douta,

        input         clkb,
        input         rstb,
        input  [8:0]  addrb,
        output [31:0] doutb
    );

    reg  [31:0]	douta_buf;
    wire [31:0]	mdouta;

    rot_SP u_arot(
        //ports
        .clka  		( clka  		),
        .rsta  		( rsta  		),
        .addra 		( addra 		),
        .douta 		( mdouta 		)
    );

    always @(posedge clka or posedge rsta) begin
        if(rsta) begin
            douta_buf <= 0;
        end
        else begin
            douta_buf <= mdouta;
        end
    end
    assign douta = douta_buf;

    reg  [31:0]	doutb_buf;
    wire [31:0]	mdoutb;

    rot_SP u_brot(
        //ports
        .clka  		( clkb  		),
        .rsta  		( rstb  		),
        .addra 		( addrb 		),
        .douta 		( mdoutb 		)
    );

    always @(posedge clkb or posedge rstb) begin
        if(rstb) begin
            doutb_buf <= 0;
        end
        else begin
            doutb_buf <= mdoutb;
        end
    end
    assign doutb = doutb_buf;

endmodule

module rot_SP (
        input         clka,
        input         rsta,
        input  [8:0]  addra,
        output [31:0] douta
    );

    reg [31:0] douta_buf;
    always @(posedge clka) begin
        if (rsta) begin
            douta_buf <= 0;
        end
        else begin
            case (addra)
                9'h0000: douta_buf <= 32'h00001000000000000000000000000000;
                9'h0001: douta_buf <= 32'h00001000000000000000000000000100;
                9'h0002: douta_buf <= 32'h00001000000000000000000000001000;
                9'h0003: douta_buf <= 32'h00001000000000000000000000001100;
                9'h0004: douta_buf <= 32'h00001000000000000000000000010000;
                9'h0005: douta_buf <= 32'h00001000000000000000000000010100;
                9'h0006: douta_buf <= 32'h00001000000000000000000000011000;
                9'h0007: douta_buf <= 32'h00001000000000000000000000011100;
                9'h0008: douta_buf <= 32'h00001000000000000000000000100000;
                9'h0009: douta_buf <= 32'h00001000000000000000000000100100;
                9'h000a: douta_buf <= 32'h00001000000000000000000000101000;
                9'h000b: douta_buf <= 32'h00001000000000000000000000101100;
                9'h000c: douta_buf <= 32'h00000111111111110000000000110000;
                9'h000d: douta_buf <= 32'h00000111111111110000000000110100;
                9'h000e: douta_buf <= 32'h00000111111111110000000000111000;
                9'h000f: douta_buf <= 32'h00000111111111110000000000111100;
                9'h0010: douta_buf <= 32'h00000111111111110000000001000000;
                9'h0011: douta_buf <= 32'h00000111111111110000000001000100;
                9'h0012: douta_buf <= 32'h00000111111111110000000001001000;
                9'h0013: douta_buf <= 32'h00000111111111110000000001001100;
                9'h0014: douta_buf <= 32'h00000111111111100000000001010000;
                9'h0015: douta_buf <= 32'h00000111111111100000000001010100;
                9'h0016: douta_buf <= 32'h00000111111111100000000001011000;
                9'h0017: douta_buf <= 32'h00000111111111100000000001011100;
                9'h0018: douta_buf <= 32'h00000111111111100000000001100000;
                9'h0019: douta_buf <= 32'h00000111111111100000000001100100;
                9'h001a: douta_buf <= 32'h00000111111111010000000001101000;
                9'h001b: douta_buf <= 32'h00000111111111010000000001101100;
                9'h001c: douta_buf <= 32'h00000111111111010000000001110000;
                9'h001d: douta_buf <= 32'h00000111111111010000000001110100;
                9'h001e: douta_buf <= 32'h00000111111111000000000001111000;
                9'h001f: douta_buf <= 32'h00000111111111000000000001111100;
                9'h0020: douta_buf <= 32'h00000111111111000000000010000000;
                9'h0021: douta_buf <= 32'h00000111111111000000000010000100;
                9'h0022: douta_buf <= 32'h00000111111110110000000010001000;
                9'h0023: douta_buf <= 32'h00000111111110110000000010001100;
                9'h0024: douta_buf <= 32'h00000111111110110000000010010000;
                9'h0025: douta_buf <= 32'h00000111111110110000000010010100;
                9'h0026: douta_buf <= 32'h00000111111110100000000010011000;
                9'h0027: douta_buf <= 32'h00000111111110100000000010011100;
                9'h0028: douta_buf <= 32'h00000111111110100000000010100000;
                9'h0029: douta_buf <= 32'h00000111111110010000000010100100;
                9'h002a: douta_buf <= 32'h00000111111110010000000010101000;
                9'h002b: douta_buf <= 32'h00000111111110010000000010101100;
                9'h002c: douta_buf <= 32'h00000111111110000000000010110000;
                9'h002d: douta_buf <= 32'h00000111111110000000000010110100;
                9'h002e: douta_buf <= 32'h00000111111110000000000010111000;
                9'h002f: douta_buf <= 32'h00000111111101110000000010111100;
                9'h0030: douta_buf <= 32'h00000111111101110000000011000000;
                9'h0031: douta_buf <= 32'h00000111111101110000000011000100;
                9'h0032: douta_buf <= 32'h00000111111101100000000011001000;
                9'h0033: douta_buf <= 32'h00000111111101100000000011001100;
                9'h0034: douta_buf <= 32'h00000111111101010000000011010000;
                9'h0035: douta_buf <= 32'h00000111111101010000000011010100;
                9'h0036: douta_buf <= 32'h00000111111101010000000011011000;
                9'h0037: douta_buf <= 32'h00000111111101000000000011011100;
                9'h0038: douta_buf <= 32'h00000111111101000000000011100000;
                9'h0039: douta_buf <= 32'h00000111111100110000000011100100;
                9'h003a: douta_buf <= 32'h00000111111100110000000011101000;
                9'h003b: douta_buf <= 32'h00000111111100100000000011101100;
                9'h003c: douta_buf <= 32'h00000111111100100000000011110000;
                9'h003d: douta_buf <= 32'h00000111111100010000000011110011;
                9'h003e: douta_buf <= 32'h00000111111100010000000011110111;
                9'h003f: douta_buf <= 32'h00000111111100010000000011111011;
                9'h0040: douta_buf <= 32'h00000111111100000000000011111111;
                9'h0041: douta_buf <= 32'h00000111111100000000000100000011;
                9'h0042: douta_buf <= 32'h00000111111011110000000100000111;
                9'h0043: douta_buf <= 32'h00000111111011100000000100001011;
                9'h0044: douta_buf <= 32'h00000111111011100000000100001111;
                9'h0045: douta_buf <= 32'h00000111111011010000000100010011;
                9'h0046: douta_buf <= 32'h00000111111011010000000100010111;
                9'h0047: douta_buf <= 32'h00000111111011000000000100011011;
                9'h0048: douta_buf <= 32'h00000111111011000000000100011111;
                9'h0049: douta_buf <= 32'h00000111111010110000000100100011;
                9'h004a: douta_buf <= 32'h00000111111010110000000100100111;
                9'h004b: douta_buf <= 32'h00000111111010100000000100101011;
                9'h004c: douta_buf <= 32'h00000111111010010000000100101111;
                9'h004d: douta_buf <= 32'h00000111111010010000000100110011;
                9'h004e: douta_buf <= 32'h00000111111010000000000100110111;
                9'h004f: douta_buf <= 32'h00000111111010000000000100111011;
                9'h0050: douta_buf <= 32'h00000111111001110000000100111111;
                9'h0051: douta_buf <= 32'h00000111111001100000000101000011;
                9'h0052: douta_buf <= 32'h00000111111001100000000101000111;
                9'h0053: douta_buf <= 32'h00000111111001010000000101001011;
                9'h0054: douta_buf <= 32'h00000111111001000000000101001111;
                9'h0055: douta_buf <= 32'h00000111111001000000000101010011;
                9'h0056: douta_buf <= 32'h00000111111000110000000101010110;
                9'h0057: douta_buf <= 32'h00000111111000100000000101011010;
                9'h0058: douta_buf <= 32'h00000111111000100000000101011110;
                9'h0059: douta_buf <= 32'h00000111111000010000000101100010;
                9'h005a: douta_buf <= 32'h00000111111000000000000101100110;
                9'h005b: douta_buf <= 32'h00000111111000000000000101101010;
                9'h005c: douta_buf <= 32'h00000111110111110000000101101110;
                9'h005d: douta_buf <= 32'h00000111110111100000000101110010;
                9'h005e: douta_buf <= 32'h00000111110111100000000101110110;
                9'h005f: douta_buf <= 32'h00000111110111010000000101111010;
                9'h0060: douta_buf <= 32'h00000111110111000000000101111110;
                9'h0061: douta_buf <= 32'h00000111110110110000000110000010;
                9'h0062: douta_buf <= 32'h00000111110110110000000110000110;
                9'h0063: douta_buf <= 32'h00000111110110100000000110001010;
                9'h0064: douta_buf <= 32'h00000111110110010000000110001110;
                9'h0065: douta_buf <= 32'h00000111110110000000000110010010;
                9'h0066: douta_buf <= 32'h00000111110101110000000110010101;
                9'h0067: douta_buf <= 32'h00000111110101110000000110011001;
                9'h0068: douta_buf <= 32'h00000111110101100000000110011101;
                9'h0069: douta_buf <= 32'h00000111110101010000000110100001;
                9'h006a: douta_buf <= 32'h00000111110101000000000110100101;
                9'h006b: douta_buf <= 32'h00000111110100110000000110101001;
                9'h006c: douta_buf <= 32'h00000111110100110000000110101101;
                9'h006d: douta_buf <= 32'h00000111110100100000000110110001;
                9'h006e: douta_buf <= 32'h00000111110100010000000110110101;
                9'h006f: douta_buf <= 32'h00000111110100000000000110111001;
                9'h0070: douta_buf <= 32'h00000111110011110000000110111101;
                9'h0071: douta_buf <= 32'h00000111110011100000000111000000;
                9'h0072: douta_buf <= 32'h00000111110011010000000111000100;
                9'h0073: douta_buf <= 32'h00000111110011010000000111001000;
                9'h0074: douta_buf <= 32'h00000111110011000000000111001100;
                9'h0075: douta_buf <= 32'h00000111110010110000000111010000;
                9'h0076: douta_buf <= 32'h00000111110010100000000111010100;
                9'h0077: douta_buf <= 32'h00000111110010010000000111011000;
                9'h0078: douta_buf <= 32'h00000111110010000000000111011100;
                9'h0079: douta_buf <= 32'h00000111110001110000000111100000;
                9'h007a: douta_buf <= 32'h00000111110001100000000111100100;
                9'h007b: douta_buf <= 32'h00000111110001010000000111100111;
                9'h007c: douta_buf <= 32'h00000111110001000000000111101011;
                9'h007d: douta_buf <= 32'h00000111110000110000000111101111;
                9'h007e: douta_buf <= 32'h00000111110000100000000111110011;
                9'h007f: douta_buf <= 32'h00000111110000010000000111110111;
                9'h0080: douta_buf <= 32'h00000111110000000000000111111011;
                9'h0081: douta_buf <= 32'h00000111101111110000000111111111;
                9'h0082: douta_buf <= 32'h00000111101111100000001000000011;
                9'h0083: douta_buf <= 32'h00000111101111010000001000000110;
                9'h0084: douta_buf <= 32'h00000111101111000000001000001010;
                9'h0085: douta_buf <= 32'h00000111101110110000001000001110;
                9'h0086: douta_buf <= 32'h00000111101110100000001000010010;
                9'h0087: douta_buf <= 32'h00000111101110010000001000010110;
                9'h0088: douta_buf <= 32'h00000111101110000000001000011010;
                9'h0089: douta_buf <= 32'h00000111101101110000001000011110;
                9'h008a: douta_buf <= 32'h00000111101101100000001000100010;
                9'h008b: douta_buf <= 32'h00000111101101010000001000100101;
                9'h008c: douta_buf <= 32'h00000111101101000000001000101001;
                9'h008d: douta_buf <= 32'h00000111101100110000001000101101;
                9'h008e: douta_buf <= 32'h00000111101100100000001000110001;
                9'h008f: douta_buf <= 32'h00000111101100010000001000110101;
                9'h0090: douta_buf <= 32'h00000111101011110000001000111001;
                9'h0091: douta_buf <= 32'h00000111101011100000001000111100;
                9'h0092: douta_buf <= 32'h00000111101011010000001001000000;
                9'h0093: douta_buf <= 32'h00000111101011000000001001000100;
                9'h0094: douta_buf <= 32'h00000111101010110000001001001000;
                9'h0095: douta_buf <= 32'h00000111101010100000001001001100;
                9'h0096: douta_buf <= 32'h00000111101010010000001001010000;
                9'h0097: douta_buf <= 32'h00000111101010000000001001010011;
                9'h0098: douta_buf <= 32'h00000111101001100000001001010111;
                9'h0099: douta_buf <= 32'h00000111101001010000001001011011;
                9'h009a: douta_buf <= 32'h00000111101001000000001001011111;
                9'h009b: douta_buf <= 32'h00000111101000110000001001100011;
                9'h009c: douta_buf <= 32'h00000111101000100000001001100111;
                9'h009d: douta_buf <= 32'h00000111101000000000001001101010;
                9'h009e: douta_buf <= 32'h00000111100111110000001001101110;
                9'h009f: douta_buf <= 32'h00000111100111100000001001110010;
                9'h00a0: douta_buf <= 32'h00000111100111010000001001110110;
                9'h00a1: douta_buf <= 32'h00000111100111000000001001111010;
                9'h00a2: douta_buf <= 32'h00000111100110100000001001111101;
                9'h00a3: douta_buf <= 32'h00000111100110010000001010000001;
                9'h00a4: douta_buf <= 32'h00000111100110000000001010000101;
                9'h00a5: douta_buf <= 32'h00000111100101110000001010001001;
                9'h00a6: douta_buf <= 32'h00000111100101010000001010001101;
                9'h00a7: douta_buf <= 32'h00000111100101000000001010010000;
                9'h00a8: douta_buf <= 32'h00000111100100110000001010010100;
                9'h00a9: douta_buf <= 32'h00000111100100010000001010011000;
                9'h00aa: douta_buf <= 32'h00000111100100000000001010011100;
                9'h00ab: douta_buf <= 32'h00000111100011110000001010100000;
                9'h00ac: douta_buf <= 32'h00000111100011010000001010100011;
                9'h00ad: douta_buf <= 32'h00000111100011000000001010100111;
                9'h00ae: douta_buf <= 32'h00000111100010110000001010101011;
                9'h00af: douta_buf <= 32'h00000111100010010000001010101111;
                9'h00b0: douta_buf <= 32'h00000111100010000000001010110010;
                9'h00b1: douta_buf <= 32'h00000111100001110000001010110110;
                9'h00b2: douta_buf <= 32'h00000111100001010000001010111010;
                9'h00b3: douta_buf <= 32'h00000111100001000000001010111110;
                9'h00b4: douta_buf <= 32'h00000111100000110000001011000001;
                9'h00b5: douta_buf <= 32'h00000111100000010000001011000101;
                9'h00b6: douta_buf <= 32'h00000111100000000000001011001001;
                9'h00b7: douta_buf <= 32'h00000111011111100000001011001101;
                9'h00b8: douta_buf <= 32'h00000111011111010000001011010000;
                9'h00b9: douta_buf <= 32'h00000111011111000000001011010100;
                9'h00ba: douta_buf <= 32'h00000111011110100000001011011000;
                9'h00bb: douta_buf <= 32'h00000111011110010000001011011100;
                9'h00bc: douta_buf <= 32'h00000111011101110000001011011111;
                9'h00bd: douta_buf <= 32'h00000111011101100000001011100011;
                9'h00be: douta_buf <= 32'h00000111011101010000001011100111;
                9'h00bf: douta_buf <= 32'h00000111011100110000001011101011;
                9'h00c0: douta_buf <= 32'h00000111011100100000001011101110;
                9'h00c1: douta_buf <= 32'h00000111011100000000001011110010;
                9'h00c2: douta_buf <= 32'h00000111011011110000001011110110;
                9'h00c3: douta_buf <= 32'h00000111011011010000001011111010;
                9'h00c4: douta_buf <= 32'h00000111011011000000001011111101;
                9'h00c5: douta_buf <= 32'h00000111011010100000001100000001;
                9'h00c6: douta_buf <= 32'h00000111011010010000001100000101;
                9'h00c7: douta_buf <= 32'h00000111011001110000001100001000;
                9'h00c8: douta_buf <= 32'h00000111011001100000001100001100;
                9'h00c9: douta_buf <= 32'h00000111011001000000001100010000;
                9'h00ca: douta_buf <= 32'h00000111011000110000001100010011;
                9'h00cb: douta_buf <= 32'h00000111011000010000001100010111;
                9'h00cc: douta_buf <= 32'h00000111010111110000001100011011;
                9'h00cd: douta_buf <= 32'h00000111010111100000001100011110;
                9'h00ce: douta_buf <= 32'h00000111010111000000001100100010;
                9'h00cf: douta_buf <= 32'h00000111010110110000001100100110;
                9'h00d0: douta_buf <= 32'h00000111010110010000001100101010;
                9'h00d1: douta_buf <= 32'h00000111010110000000001100101101;
                9'h00d2: douta_buf <= 32'h00000111010101100000001100110001;
                9'h00d3: douta_buf <= 32'h00000111010101000000001100110101;
                9'h00d4: douta_buf <= 32'h00000111010100110000001100111000;
                9'h00d5: douta_buf <= 32'h00000111010100010000001100111100;
                9'h00d6: douta_buf <= 32'h00000111010100000000001101000000;
                9'h00d7: douta_buf <= 32'h00000111010011100000001101000011;
                9'h00d8: douta_buf <= 32'h00000111010011000000001101000111;
                9'h00d9: douta_buf <= 32'h00000111010010110000001101001010;
                9'h00da: douta_buf <= 32'h00000111010010010000001101001110;
                9'h00db: douta_buf <= 32'h00000111010001110000001101010010;
                9'h00dc: douta_buf <= 32'h00000111010001100000001101010101;
                9'h00dd: douta_buf <= 32'h00000111010001000000001101011001;
                9'h00de: douta_buf <= 32'h00000111010000100000001101011101;
                9'h00df: douta_buf <= 32'h00000111010000010000001101100000;
                9'h00e0: douta_buf <= 32'h00000111001111110000001101100100;
                9'h00e1: douta_buf <= 32'h00000111001111010000001101101000;
                9'h00e2: douta_buf <= 32'h00000111001111000000001101101011;
                9'h00e3: douta_buf <= 32'h00000111001110100000001101101111;
                9'h00e4: douta_buf <= 32'h00000111001110000000001101110010;
                9'h00e5: douta_buf <= 32'h00000111001101100000001101110110;
                9'h00e6: douta_buf <= 32'h00000111001101010000001101111010;
                9'h00e7: douta_buf <= 32'h00000111001100110000001101111101;
                9'h00e8: douta_buf <= 32'h00000111001100010000001110000001;
                9'h00e9: douta_buf <= 32'h00000111001011110000001110000100;
                9'h00ea: douta_buf <= 32'h00000111001011100000001110001000;
                9'h00eb: douta_buf <= 32'h00000111001011000000001110001100;
                9'h00ec: douta_buf <= 32'h00000111001010100000001110001111;
                9'h00ed: douta_buf <= 32'h00000111001010000000001110010011;
                9'h00ee: douta_buf <= 32'h00000111001001110000001110010110;
                9'h00ef: douta_buf <= 32'h00000111001001010000001110011010;
                9'h00f0: douta_buf <= 32'h00000111001000110000001110011101;
                9'h00f1: douta_buf <= 32'h00000111001000010000001110100001;
                9'h00f2: douta_buf <= 32'h00000111000111110000001110100101;
                9'h00f3: douta_buf <= 32'h00000111000111100000001110101000;
                9'h00f4: douta_buf <= 32'h00000111000111000000001110101100;
                9'h00f5: douta_buf <= 32'h00000111000110100000001110101111;
                9'h00f6: douta_buf <= 32'h00000111000110000000001110110011;
                9'h00f7: douta_buf <= 32'h00000111000101100000001110110110;
                9'h00f8: douta_buf <= 32'h00000111000101000000001110111010;
                9'h00f9: douta_buf <= 32'h00000111000100100000001110111101;
                9'h00fa: douta_buf <= 32'h00000111000100010000001111000001;
                9'h00fb: douta_buf <= 32'h00000111000011110000001111000101;
                9'h00fc: douta_buf <= 32'h00000111000011010000001111001000;
                9'h00fd: douta_buf <= 32'h00000111000010110000001111001100;
                9'h00fe: douta_buf <= 32'h00000111000010010000001111001111;
                9'h00ff: douta_buf <= 32'h00000111000001110000001111010011;
                9'h0100: douta_buf <= 32'h00000111000001010000001111010110;
                9'h0101: douta_buf <= 32'h00000111000000110000001111011010;
                9'h0102: douta_buf <= 32'h00000111000000010000001111011101;
                9'h0103: douta_buf <= 32'h00000110111111110000001111100001;
                9'h0104: douta_buf <= 32'h00000110111111010000001111100100;
                9'h0105: douta_buf <= 32'h00000110111110110000001111101000;
                9'h0106: douta_buf <= 32'h00000110111110100000001111101011;
                9'h0107: douta_buf <= 32'h00000110111110000000001111101111;
                9'h0108: douta_buf <= 32'h00000110111101100000001111110010;
                9'h0109: douta_buf <= 32'h00000110111101000000001111110110;
                9'h010a: douta_buf <= 32'h00000110111100100000001111111001;
                9'h010b: douta_buf <= 32'h00000110111100000000001111111101;
                9'h010c: douta_buf <= 32'h00000110111011100000010000000000;
                9'h010d: douta_buf <= 32'h00000110111011000000010000000011;
                9'h010e: douta_buf <= 32'h00000110111010100000010000000111;
                9'h010f: douta_buf <= 32'h00000110111010000000010000001010;
                9'h0110: douta_buf <= 32'h00000110111001100000010000001110;
                9'h0111: douta_buf <= 32'h00000110111001000000010000010001;
                9'h0112: douta_buf <= 32'h00000110111000010000010000010101;
                9'h0113: douta_buf <= 32'h00000110110111110000010000011000;
                9'h0114: douta_buf <= 32'h00000110110111010000010000011100;
                9'h0115: douta_buf <= 32'h00000110110110110000010000011111;
                9'h0116: douta_buf <= 32'h00000110110110010000010000100010;
                9'h0117: douta_buf <= 32'h00000110110101110000010000100110;
                9'h0118: douta_buf <= 32'h00000110110101010000010000101001;
                9'h0119: douta_buf <= 32'h00000110110100110000010000101101;
                9'h011a: douta_buf <= 32'h00000110110100010000010000110000;
                9'h011b: douta_buf <= 32'h00000110110011110000010000110100;
                9'h011c: douta_buf <= 32'h00000110110011010000010000110111;
                9'h011d: douta_buf <= 32'h00000110110010110000010000111010;
                9'h011e: douta_buf <= 32'h00000110110010010000010000111110;
                9'h011f: douta_buf <= 32'h00000110110001100000010001000001;
                9'h0120: douta_buf <= 32'h00000110110001000000010001000101;
                9'h0121: douta_buf <= 32'h00000110110000100000010001001000;
                9'h0122: douta_buf <= 32'h00000110110000000000010001001011;
                9'h0123: douta_buf <= 32'h00000110101111100000010001001111;
                9'h0124: douta_buf <= 32'h00000110101111000000010001010010;
                9'h0125: douta_buf <= 32'h00000110101110100000010001010101;
                9'h0126: douta_buf <= 32'h00000110101101110000010001011001;
                9'h0127: douta_buf <= 32'h00000110101101010000010001011100;
                9'h0128: douta_buf <= 32'h00000110101100110000010001011111;
                9'h0129: douta_buf <= 32'h00000110101100010000010001100011;
                9'h012a: douta_buf <= 32'h00000110101011110000010001100110;
                9'h012b: douta_buf <= 32'h00000110101011000000010001101001;
                9'h012c: douta_buf <= 32'h00000110101010100000010001101101;
                9'h012d: douta_buf <= 32'h00000110101010000000010001110000;
                9'h012e: douta_buf <= 32'h00000110101001100000010001110011;
                9'h012f: douta_buf <= 32'h00000110101001000000010001110111;
                9'h0130: douta_buf <= 32'h00000110101000010000010001111010;
                9'h0131: douta_buf <= 32'h00000110100111110000010001111101;
                9'h0132: douta_buf <= 32'h00000110100111010000010010000001;
                9'h0133: douta_buf <= 32'h00000110100110110000010010000100;
                9'h0134: douta_buf <= 32'h00000110100110000000010010000111;
                9'h0135: douta_buf <= 32'h00000110100101100000010010001011;
                9'h0136: douta_buf <= 32'h00000110100101000000010010001110;
                9'h0137: douta_buf <= 32'h00000110100100010000010010010001;
                9'h0138: douta_buf <= 32'h00000110100011110000010010010100;
                9'h0139: douta_buf <= 32'h00000110100011010000010010011000;
                9'h013a: douta_buf <= 32'h00000110100010110000010010011011;
                9'h013b: douta_buf <= 32'h00000110100010000000010010011110;
                9'h013c: douta_buf <= 32'h00000110100001100000010010100010;
                9'h013d: douta_buf <= 32'h00000110100001000000010010100101;
                9'h013e: douta_buf <= 32'h00000110100000010000010010101000;
                9'h013f: douta_buf <= 32'h00000110011111110000010010101011;
                9'h0140: douta_buf <= 32'h00000110011111010000010010101111;
                9'h0141: douta_buf <= 32'h00000110011110100000010010110010;
                9'h0142: douta_buf <= 32'h00000110011110000000010010110101;
                9'h0143: douta_buf <= 32'h00000110011101100000010010111000;
                9'h0144: douta_buf <= 32'h00000110011100110000010010111100;
                9'h0145: douta_buf <= 32'h00000110011100010000010010111111;
                9'h0146: douta_buf <= 32'h00000110011011100000010011000010;
                9'h0147: douta_buf <= 32'h00000110011011000000010011000101;
                9'h0148: douta_buf <= 32'h00000110011010100000010011001000;
                9'h0149: douta_buf <= 32'h00000110011001110000010011001100;
                9'h014a: douta_buf <= 32'h00000110011001010000010011001111;
                9'h014b: douta_buf <= 32'h00000110011000100000010011010010;
                9'h014c: douta_buf <= 32'h00000110011000000000010011010101;
                9'h014d: douta_buf <= 32'h00000110010111100000010011011000;
                9'h014e: douta_buf <= 32'h00000110010110110000010011011100;
                9'h014f: douta_buf <= 32'h00000110010110010000010011011111;
                9'h0150: douta_buf <= 32'h00000110010101100000010011100010;
                9'h0151: douta_buf <= 32'h00000110010101000000010011100101;
                9'h0152: douta_buf <= 32'h00000110010100010000010011101000;
                9'h0153: douta_buf <= 32'h00000110010011110000010011101011;
                9'h0154: douta_buf <= 32'h00000110010011010000010011101111;
                9'h0155: douta_buf <= 32'h00000110010010100000010011110010;
                9'h0156: douta_buf <= 32'h00000110010010000000010011110101;
                9'h0157: douta_buf <= 32'h00000110010001010000010011111000;
                9'h0158: douta_buf <= 32'h00000110010000110000010011111011;
                9'h0159: douta_buf <= 32'h00000110010000000000010011111110;
                9'h015a: douta_buf <= 32'h00000110001111100000010100000001;
                9'h015b: douta_buf <= 32'h00000110001110110000010100000100;
                9'h015c: douta_buf <= 32'h00000110001110010000010100001000;
                9'h015d: douta_buf <= 32'h00000110001101100000010100001011;
                9'h015e: douta_buf <= 32'h00000110001101000000010100001110;
                9'h015f: douta_buf <= 32'h00000110001100010000010100010001;
                9'h0160: douta_buf <= 32'h00000110001011100000010100010100;
                9'h0161: douta_buf <= 32'h00000110001011000000010100010111;
                9'h0162: douta_buf <= 32'h00000110001010010000010100011010;
                9'h0163: douta_buf <= 32'h00000110001001110000010100011101;
                9'h0164: douta_buf <= 32'h00000110001001000000010100100000;
                9'h0165: douta_buf <= 32'h00000110001000100000010100100011;
                9'h0166: douta_buf <= 32'h00000110000111110000010100100110;
                9'h0167: douta_buf <= 32'h00000110000111010000010100101010;
                9'h0168: douta_buf <= 32'h00000110000110100000010100101101;
                9'h0169: douta_buf <= 32'h00000110000101110000010100110000;
                9'h016a: douta_buf <= 32'h00000110000101010000010100110011;
                9'h016b: douta_buf <= 32'h00000110000100100000010100110110;
                9'h016c: douta_buf <= 32'h00000110000100000000010100111001;
                9'h016d: douta_buf <= 32'h00000110000011010000010100111100;
                9'h016e: douta_buf <= 32'h00000110000010100000010100111111;
                9'h016f: douta_buf <= 32'h00000110000010000000010101000010;
                9'h0170: douta_buf <= 32'h00000110000001010000010101000101;
                9'h0171: douta_buf <= 32'h00000110000000100000010101001000;
                9'h0172: douta_buf <= 32'h00000110000000000000010101001011;
                9'h0173: douta_buf <= 32'h00000101111111010000010101001110;
                9'h0174: douta_buf <= 32'h00000101111110100000010101010001;
                9'h0175: douta_buf <= 32'h00000101111110000000010101010100;
                9'h0176: douta_buf <= 32'h00000101111101010000010101010111;
                9'h0177: douta_buf <= 32'h00000101111100100000010101011010;
                9'h0178: douta_buf <= 32'h00000101111100000000010101011101;
                9'h0179: douta_buf <= 32'h00000101111011010000010101100000;
                9'h017a: douta_buf <= 32'h00000101111010100000010101100011;
                9'h017b: douta_buf <= 32'h00000101111010000000010101100110;
                9'h017c: douta_buf <= 32'h00000101111001010000010101101001;
                9'h017d: douta_buf <= 32'h00000101111000100000010101101100;
                9'h017e: douta_buf <= 32'h00000101111000000000010101101110;
                9'h017f: douta_buf <= 32'h00000101110111010000010101110001;
                9'h0180: douta_buf <= 32'h00000101110110100000010101110100;
                9'h0181: douta_buf <= 32'h00000101110101110000010101110111;
                9'h0182: douta_buf <= 32'h00000101110101010000010101111010;
                9'h0183: douta_buf <= 32'h00000101110100100000010101111101;
                9'h0184: douta_buf <= 32'h00000101110011110000010110000000;
                9'h0185: douta_buf <= 32'h00000101110011000000010110000011;
                9'h0186: douta_buf <= 32'h00000101110010100000010110000110;
                9'h0187: douta_buf <= 32'h00000101110001110000010110001001;
                9'h0188: douta_buf <= 32'h00000101110001000000010110001100;
                9'h0189: douta_buf <= 32'h00000101110000010000010110001110;
                9'h018a: douta_buf <= 32'h00000101101111110000010110010001;
                9'h018b: douta_buf <= 32'h00000101101111000000010110010100;
                9'h018c: douta_buf <= 32'h00000101101110010000010110010111;
                9'h018d: douta_buf <= 32'h00000101101101100000010110011010;
                9'h018e: douta_buf <= 32'h00000101101100110000010110011101;
                9'h018f: douta_buf <= 32'h00000101101100010000010110100000;
                9'h0190: douta_buf <= 32'h00000101101011100000010110100010;
                9'h0191: douta_buf <= 32'h00000101101010110000010110100101;
                9'h0192: douta_buf <= 32'h00000101101010000000010110101000;
                9'h0193: douta_buf <= 32'h00000101101001010000010110101011;
                9'h0194: douta_buf <= 32'h00000101101000100000010110101110;
                9'h0195: douta_buf <= 32'h00000101101000000000010110110001;
                9'h0196: douta_buf <= 32'h00000101100111010000010110110011;
                9'h0197: douta_buf <= 32'h00000101100110100000010110110110;
                9'h0198: douta_buf <= 32'h00000101100101110000010110111001;
                9'h0199: douta_buf <= 32'h00000101100101000000010110111100;
                9'h019a: douta_buf <= 32'h00000101100100010000010110111111;
                9'h019b: douta_buf <= 32'h00000101100011100000010111000001;
                9'h019c: douta_buf <= 32'h00000101100011000000010111000100;
                9'h019d: douta_buf <= 32'h00000101100010010000010111000111;
                9'h019e: douta_buf <= 32'h00000101100001100000010111001010;
                9'h019f: douta_buf <= 32'h00000101100000110000010111001100;
                9'h01a0: douta_buf <= 32'h00000101100000000000010111001111;
                9'h01a1: douta_buf <= 32'h00000101011111010000010111010010;
                9'h01a2: douta_buf <= 32'h00000101011110100000010111010101;
                9'h01a3: douta_buf <= 32'h00000101011101110000010111010111;
                9'h01a4: douta_buf <= 32'h00000101011101000000010111011010;
                9'h01a5: douta_buf <= 32'h00000101011100010000010111011101;
                9'h01a6: douta_buf <= 32'h00000101011011100000010111100000;
                9'h01a7: douta_buf <= 32'h00000101011011000000010111100010;
                9'h01a8: douta_buf <= 32'h00000101011010010000010111100101;
                9'h01a9: douta_buf <= 32'h00000101011001100000010111101000;
                9'h01aa: douta_buf <= 32'h00000101011000110000010111101010;
                9'h01ab: douta_buf <= 32'h00000101011000000000010111101101;
                9'h01ac: douta_buf <= 32'h00000101010111010000010111110000;
                9'h01ad: douta_buf <= 32'h00000101010110100000010111110010;
                9'h01ae: douta_buf <= 32'h00000101010101110000010111110101;
                9'h01af: douta_buf <= 32'h00000101010101000000010111111000;
                9'h01b0: douta_buf <= 32'h00000101010100010000010111111010;
                9'h01b1: douta_buf <= 32'h00000101010011100000010111111101;
                9'h01b2: douta_buf <= 32'h00000101010010110000011000000000;
                9'h01b3: douta_buf <= 32'h00000101010010000000011000000010;
                9'h01b4: douta_buf <= 32'h00000101010001010000011000000101;
                9'h01b5: douta_buf <= 32'h00000101010000100000011000001000;
                9'h01b6: douta_buf <= 32'h00000101001111110000011000001010;
                9'h01b7: douta_buf <= 32'h00000101001111000000011000001101;
                9'h01b8: douta_buf <= 32'h00000101001110010000011000010000;
                9'h01b9: douta_buf <= 32'h00000101001101100000011000010010;
                9'h01ba: douta_buf <= 32'h00000101001100110000011000010101;
                9'h01bb: douta_buf <= 32'h00000101001100000000011000010111;
                9'h01bc: douta_buf <= 32'h00000101001011010000011000011010;
                9'h01bd: douta_buf <= 32'h00000101001010100000011000011101;
                9'h01be: douta_buf <= 32'h00000101001001100000011000011111;
                9'h01bf: douta_buf <= 32'h00000101001000110000011000100010;
                9'h01c0: douta_buf <= 32'h00000101001000000000011000100100;
                9'h01c1: douta_buf <= 32'h00000101000111010000011000100111;
                9'h01c2: douta_buf <= 32'h00000101000110100000011000101001;
                9'h01c3: douta_buf <= 32'h00000101000101110000011000101100;
                9'h01c4: douta_buf <= 32'h00000101000101000000011000101110;
                9'h01c5: douta_buf <= 32'h00000101000100010000011000110001;
                9'h01c6: douta_buf <= 32'h00000101000011100000011000110100;
                9'h01c7: douta_buf <= 32'h00000101000010110000011000110110;
                9'h01c8: douta_buf <= 32'h00000101000010000000011000111001;
                9'h01c9: douta_buf <= 32'h00000101000001000000011000111011;
                9'h01ca: douta_buf <= 32'h00000101000000010000011000111110;
                9'h01cb: douta_buf <= 32'h00000100111111100000011001000000;
                9'h01cc: douta_buf <= 32'h00000100111110110000011001000011;
                9'h01cd: douta_buf <= 32'h00000100111110000000011001000101;
                9'h01ce: douta_buf <= 32'h00000100111101010000011001001000;
                9'h01cf: douta_buf <= 32'h00000100111100100000011001001010;
                9'h01d0: douta_buf <= 32'h00000100111011110000011001001101;
                9'h01d1: douta_buf <= 32'h00000100111010110000011001001111;
                9'h01d2: douta_buf <= 32'h00000100111010000000011001010001;
                9'h01d3: douta_buf <= 32'h00000100111001010000011001010100;
                9'h01d4: douta_buf <= 32'h00000100111000100000011001010110;
                9'h01d5: douta_buf <= 32'h00000100110111110000011001011001;
                9'h01d6: douta_buf <= 32'h00000100110111000000011001011011;
                9'h01d7: douta_buf <= 32'h00000100110110000000011001011110;
                9'h01d8: douta_buf <= 32'h00000100110101010000011001100000;
                9'h01d9: douta_buf <= 32'h00000100110100100000011001100010;
                9'h01da: douta_buf <= 32'h00000100110011110000011001100101;
                9'h01db: douta_buf <= 32'h00000100110011000000011001100111;
                9'h01dc: douta_buf <= 32'h00000100110010000000011001101010;
                9'h01dd: douta_buf <= 32'h00000100110001010000011001101100;
                9'h01de: douta_buf <= 32'h00000100110000100000011001101110;
                9'h01df: douta_buf <= 32'h00000100101111110000011001110001;
                9'h01e0: douta_buf <= 32'h00000100101111000000011001110011;
                9'h01e1: douta_buf <= 32'h00000100101110000000011001110110;
                9'h01e2: douta_buf <= 32'h00000100101101010000011001111000;
                9'h01e3: douta_buf <= 32'h00000100101100100000011001111010;
                9'h01e4: douta_buf <= 32'h00000100101011110000011001111101;
                9'h01e5: douta_buf <= 32'h00000100101010110000011001111111;
                9'h01e6: douta_buf <= 32'h00000100101010000000011010000001;
                9'h01e7: douta_buf <= 32'h00000100101001010000011010000100;
                9'h01e8: douta_buf <= 32'h00000100101000100000011010000110;
                9'h01e9: douta_buf <= 32'h00000100100111100000011010001000;
                9'h01ea: douta_buf <= 32'h00000100100110110000011010001011;
                9'h01eb: douta_buf <= 32'h00000100100110000000011010001101;
                9'h01ec: douta_buf <= 32'h00000100100101000000011010001111;
                9'h01ed: douta_buf <= 32'h00000100100100010000011010010001;
                9'h01ee: douta_buf <= 32'h00000100100011100000011010010100;
                9'h01ef: douta_buf <= 32'h00000100100010110000011010010110;
                9'h01f0: douta_buf <= 32'h00000100100001110000011010011000;
                9'h01f1: douta_buf <= 32'h00000100100001000000011010011011;
                9'h01f2: douta_buf <= 32'h00000100100000010000011010011101;
                9'h01f3: douta_buf <= 32'h00000100011111010000011010011111;
                9'h01f4: douta_buf <= 32'h00000100011110100000011010100001;
                9'h01f5: douta_buf <= 32'h00000100011101110000011010100100;
                9'h01f6: douta_buf <= 32'h00000100011100110000011010100110;
                9'h01f7: douta_buf <= 32'h00000100011100000000011010101000;
                9'h01f8: douta_buf <= 32'h00000100011011010000011010101010;
                9'h01f9: douta_buf <= 32'h00000100011010010000011010101100;
                9'h01fa: douta_buf <= 32'h00000100011001100000011010101111;
                9'h01fb: douta_buf <= 32'h00000100011000110000011010110001;
                9'h01fc: douta_buf <= 32'h00000100010111110000011010110011;
                9'h01fd: douta_buf <= 32'h00000100010111000000011010110101;
                9'h01fe: douta_buf <= 32'h00000100010110010000011010110111;
                9'h01ff: douta_buf <= 32'h00000100010101010000011010111010;
            endcase
        end
    end

    assign douta = douta_buf;
endmodule
module deinter (
        input         clka,
        input         rsta,
        input  [11:0] addra,
        output [21:0] douta
    );

    reg [21:0] douta_buf;
    always @(posedge clka) begin
        if (rsta) begin
            douta_buf <= 0;
        end
        else begin
            case (addra)
                12'h0000: douta_buf <= 22'h0000000000000000000000;
                12'h0001: douta_buf <= 22'h0000000000000000000000;
                12'h0002: douta_buf <= 22'h0000000000000000000000;
                12'h0003: douta_buf <= 22'h0000000000000000000000;
                12'h0004: douta_buf <= 22'h0000000000000000000000;
                12'h0005: douta_buf <= 22'h0000000000000000000000;
                12'h0006: douta_buf <= 22'h0000000000000000000000;
                12'h0007: douta_buf <= 22'h0000000000000000000000;
                12'h0008: douta_buf <= 22'h0000000000000111100010;
                12'h0009: douta_buf <= 22'h0000000000000011101000;
                12'h000a: douta_buf <= 22'h0000000000000001100110;
                12'h000b: douta_buf <= 22'h0000000000000000100000;
                12'h000c: douta_buf <= 22'h0000000000001010100111;
                12'h000d: douta_buf <= 22'h0000000000000101001101;
                12'h000e: douta_buf <= 22'h0000000000000010011011;
                12'h000f: douta_buf <= 22'h0000000000000000111101;
                12'h0010: douta_buf <= 22'h0000000000001110000100;
                12'h0011: douta_buf <= 22'h0000000000001110100011;
                12'h0012: douta_buf <= 22'h0000000000001111011100;
                12'h0013: douta_buf <= 22'h0000000000010000101111;
                12'h0014: douta_buf <= 22'h0000000000010010011100;
                12'h0015: douta_buf <= 22'h0000000000010100111101;
                12'h0016: douta_buf <= 22'h0000000000011000010010;
                12'h0017: douta_buf <= 22'h0000000000011100000001;
                12'h0018: douta_buf <= 22'h0000000000000000000000;
                12'h0019: douta_buf <= 22'h0000000000000000000000;
                12'h001a: douta_buf <= 22'h0000000000000000000000;
                12'h001b: douta_buf <= 22'h0000000000000000000000;
                12'h001c: douta_buf <= 22'h0000000000000000000000;
                12'h001d: douta_buf <= 22'h0000000000000000000000;
                12'h001e: douta_buf <= 22'h0000000000000000000000;
                12'h001f: douta_buf <= 22'h0000000000000000000000;
                12'h0020: douta_buf <= 22'h0000000000001100000010;
                12'h0021: douta_buf <= 22'h0000011000100100000010;
                12'h0022: douta_buf <= 22'h0000110000111100000010;
                12'h0023: douta_buf <= 22'h0001001001010100000010;
                12'h0024: douta_buf <= 22'h0001100001101100000010;
                12'h0025: douta_buf <= 22'h0001111010000100000010;
                12'h0026: douta_buf <= 22'h0010010010011100000010;
                12'h0027: douta_buf <= 22'h0010101010110100000010;
                12'h0028: douta_buf <= 22'h0000000100010000000010;
                12'h0029: douta_buf <= 22'h0000011100101000000010;
                12'h002a: douta_buf <= 22'h0000110101000000000010;
                12'h002b: douta_buf <= 22'h0001001101011000000010;
                12'h002c: douta_buf <= 22'h0001100101110000000010;
                12'h002d: douta_buf <= 22'h0001111110001000000010;
                12'h002e: douta_buf <= 22'h0010010110100000000010;
                12'h002f: douta_buf <= 22'h0010101110111000000010;
                12'h0030: douta_buf <= 22'h0000001000010100000010;
                12'h0031: douta_buf <= 22'h0000100000101100000010;
                12'h0032: douta_buf <= 22'h0000111001000100000010;
                12'h0033: douta_buf <= 22'h0001010001011100000010;
                12'h0034: douta_buf <= 22'h0001101001110100000010;
                12'h0035: douta_buf <= 22'h0010000010001100000010;
                12'h0036: douta_buf <= 22'h0010011010100100000010;
                12'h0037: douta_buf <= 22'h0010110010111100000010;
                12'h0038: douta_buf <= 22'h0001100000000000000001;
                12'h0039: douta_buf <= 22'h0000000000000000000000;
                12'h003a: douta_buf <= 22'h0000000000000000000000;
                12'h003b: douta_buf <= 22'h0000000000000000000000;
                12'h003c: douta_buf <= 22'h0000000000000000000000;
                12'h003d: douta_buf <= 22'h0000000000001100000010;
                12'h003e: douta_buf <= 22'h0100011000100100000010;
                12'h003f: douta_buf <= 22'h1000011000100100000010;
                12'h0040: douta_buf <= 22'h0000110000111100000010;
                12'h0041: douta_buf <= 22'h0101001001010100000010;
                12'h0042: douta_buf <= 22'h1001001001010100000010;
                12'h0043: douta_buf <= 22'h0001100001101100000010;
                12'h0044: douta_buf <= 22'h0101111010000100000010;
                12'h0045: douta_buf <= 22'h1001111010000100000010;
                12'h0046: douta_buf <= 22'h0010010010011100000010;
                12'h0047: douta_buf <= 22'h0110101010110100000010;
                12'h0048: douta_buf <= 22'h1010101010110100000010;
                12'h0049: douta_buf <= 22'h0000000100010000000010;
                12'h004a: douta_buf <= 22'h0100011100101000000010;
                12'h004b: douta_buf <= 22'h1000011100101000000010;
                12'h004c: douta_buf <= 22'h0000110101000000000010;
                12'h004d: douta_buf <= 22'h0101001101011000000010;
                12'h004e: douta_buf <= 22'h1001001101011000000010;
                12'h004f: douta_buf <= 22'h0001100101110000000010;
                12'h0050: douta_buf <= 22'h0101111110001000000010;
                12'h0051: douta_buf <= 22'h1001111110001000000010;
                12'h0052: douta_buf <= 22'h0010010110100000000010;
                12'h0053: douta_buf <= 22'h0110101110111000000010;
                12'h0054: douta_buf <= 22'h1010101110111000000010;
                12'h0055: douta_buf <= 22'h0000001000010100000010;
                12'h0056: douta_buf <= 22'h0100100000101100000010;
                12'h0057: douta_buf <= 22'h1000100000101100000010;
                12'h0058: douta_buf <= 22'h0000111001000100000010;
                12'h0059: douta_buf <= 22'h0101010001011100000010;
                12'h005a: douta_buf <= 22'h1001010001011100000010;
                12'h005b: douta_buf <= 22'h0001101001110100000010;
                12'h005c: douta_buf <= 22'h0110000010001100000010;
                12'h005d: douta_buf <= 22'h1010000010001100000010;
                12'h005e: douta_buf <= 22'h0010011010100100000010;
                12'h005f: douta_buf <= 22'h0110110010111100000010;
                12'h0060: douta_buf <= 22'h1010110010111100000010;
                12'h0061: douta_buf <= 22'h0001100000000000000001;
                12'h0062: douta_buf <= 22'h0000000000000000000000;
                12'h0063: douta_buf <= 22'h0000000000000000000000;
                12'h0064: douta_buf <= 22'h0000000000000000000000;
                12'h0065: douta_buf <= 22'h0000000000000000000000;
                12'h0066: douta_buf <= 22'h0000000000001100000010;
                12'h0067: douta_buf <= 22'h0000011000100100000010;
                12'h0068: douta_buf <= 22'h0000110000111100000010;
                12'h0069: douta_buf <= 22'h0001001001010100000010;
                12'h006a: douta_buf <= 22'h0001100001101100000010;
                12'h006b: douta_buf <= 22'h0001111010000100000010;
                12'h006c: douta_buf <= 22'h0010010010011100000010;
                12'h006d: douta_buf <= 22'h0010101010110100000010;
                12'h006e: douta_buf <= 22'h0000000000001100100110;
                12'h006f: douta_buf <= 22'h0000011000100100100110;
                12'h0070: douta_buf <= 22'h0000110000111100100110;
                12'h0071: douta_buf <= 22'h0001001001010100100110;
                12'h0072: douta_buf <= 22'h0001100001101100100110;
                12'h0073: douta_buf <= 22'h0001111010000100100110;
                12'h0074: douta_buf <= 22'h0010010010011100100110;
                12'h0075: douta_buf <= 22'h0010101010110100100110;
                12'h0076: douta_buf <= 22'h0000000100010000000010;
                12'h0077: douta_buf <= 22'h0000011100101000000010;
                12'h0078: douta_buf <= 22'h0000110101000000000010;
                12'h0079: douta_buf <= 22'h0001001101011000000010;
                12'h007a: douta_buf <= 22'h0001100101110000000010;
                12'h007b: douta_buf <= 22'h0001111110001000000010;
                12'h007c: douta_buf <= 22'h0010010110100000000010;
                12'h007d: douta_buf <= 22'h0010101110111000000010;
                12'h007e: douta_buf <= 22'h0000000100010000100110;
                12'h007f: douta_buf <= 22'h0000011100101000100110;
                12'h0080: douta_buf <= 22'h0000110101000000100110;
                12'h0081: douta_buf <= 22'h0001001101011000100110;
                12'h0082: douta_buf <= 22'h0001100101110000100110;
                12'h0083: douta_buf <= 22'h0001111110001000100110;
                12'h0084: douta_buf <= 22'h0010010110100000100110;
                12'h0085: douta_buf <= 22'h0010101110111000100110;
                12'h0086: douta_buf <= 22'h0000001000010100000010;
                12'h0087: douta_buf <= 22'h0000100000101100000010;
                12'h0088: douta_buf <= 22'h0000111001000100000010;
                12'h0089: douta_buf <= 22'h0001010001011100000010;
                12'h008a: douta_buf <= 22'h0001101001110100000010;
                12'h008b: douta_buf <= 22'h0010000010001100000010;
                12'h008c: douta_buf <= 22'h0010011010100100000010;
                12'h008d: douta_buf <= 22'h0010110010111100000010;
                12'h008e: douta_buf <= 22'h0000001000010100100110;
                12'h008f: douta_buf <= 22'h0000100000101100100110;
                12'h0090: douta_buf <= 22'h0000111001000100100110;
                12'h0091: douta_buf <= 22'h0001010001011100100110;
                12'h0092: douta_buf <= 22'h0001101001110100100110;
                12'h0093: douta_buf <= 22'h0010000010001100100110;
                12'h0094: douta_buf <= 22'h0010011010100100100110;
                12'h0095: douta_buf <= 22'h0010110010111100100110;
                12'h0096: douta_buf <= 22'h0001100000000000000001;
                12'h0097: douta_buf <= 22'h0000000000000000000000;
                12'h0098: douta_buf <= 22'h0000000000000000000000;
                12'h0099: douta_buf <= 22'h0000000000000000000000;
                12'h009a: douta_buf <= 22'h0000000000000000000000;
                12'h009b: douta_buf <= 22'h0000000000001100000010;
                12'h009c: douta_buf <= 22'h0100011000100100000010;
                12'h009d: douta_buf <= 22'h1000011000100100000010;
                12'h009e: douta_buf <= 22'h0000110000111100000010;
                12'h009f: douta_buf <= 22'h0101001001010100000010;
                12'h00a0: douta_buf <= 22'h1001001001010100000010;
                12'h00a1: douta_buf <= 22'h0001100001101100000010;
                12'h00a2: douta_buf <= 22'h0101111010000100000010;
                12'h00a3: douta_buf <= 22'h1001111010000100000010;
                12'h00a4: douta_buf <= 22'h0010010010011100000010;
                12'h00a5: douta_buf <= 22'h0110101010110100000010;
                12'h00a6: douta_buf <= 22'h1010101010110100000010;
                12'h00a7: douta_buf <= 22'h0000000000001100100110;
                12'h00a8: douta_buf <= 22'h0100011000100100100110;
                12'h00a9: douta_buf <= 22'h1000011000100100100110;
                12'h00aa: douta_buf <= 22'h0000110000111100100110;
                12'h00ab: douta_buf <= 22'h0101001001010100100110;
                12'h00ac: douta_buf <= 22'h1001001001010100100110;
                12'h00ad: douta_buf <= 22'h0001100001101100100110;
                12'h00ae: douta_buf <= 22'h0101111010000100100110;
                12'h00af: douta_buf <= 22'h1001111010000100100110;
                12'h00b0: douta_buf <= 22'h0010010010011100100110;
                12'h00b1: douta_buf <= 22'h0110101010110100100110;
                12'h00b2: douta_buf <= 22'h1010101010110100100110;
                12'h00b3: douta_buf <= 22'h0000000100010000000010;
                12'h00b4: douta_buf <= 22'h0100011100101000000010;
                12'h00b5: douta_buf <= 22'h1000011100101000000010;
                12'h00b6: douta_buf <= 22'h0000110101000000000010;
                12'h00b7: douta_buf <= 22'h0101001101011000000010;
                12'h00b8: douta_buf <= 22'h1001001101011000000010;
                12'h00b9: douta_buf <= 22'h0001100101110000000010;
                12'h00ba: douta_buf <= 22'h0101111110001000000010;
                12'h00bb: douta_buf <= 22'h1001111110001000000010;
                12'h00bc: douta_buf <= 22'h0010010110100000000010;
                12'h00bd: douta_buf <= 22'h0110101110111000000010;
                12'h00be: douta_buf <= 22'h1010101110111000000010;
                12'h00bf: douta_buf <= 22'h0000000100010000100110;
                12'h00c0: douta_buf <= 22'h0100011100101000100110;
                12'h00c1: douta_buf <= 22'h1000011100101000100110;
                12'h00c2: douta_buf <= 22'h0000110101000000100110;
                12'h00c3: douta_buf <= 22'h0101001101011000100110;
                12'h00c4: douta_buf <= 22'h1001001101011000100110;
                12'h00c5: douta_buf <= 22'h0001100101110000100110;
                12'h00c6: douta_buf <= 22'h0101111110001000100110;
                12'h00c7: douta_buf <= 22'h1001111110001000100110;
                12'h00c8: douta_buf <= 22'h0010010110100000100110;
                12'h00c9: douta_buf <= 22'h0110101110111000100110;
                12'h00ca: douta_buf <= 22'h1010101110111000100110;
                12'h00cb: douta_buf <= 22'h0000001000010100000010;
                12'h00cc: douta_buf <= 22'h0100100000101100000010;
                12'h00cd: douta_buf <= 22'h1000100000101100000010;
                12'h00ce: douta_buf <= 22'h0000111001000100000010;
                12'h00cf: douta_buf <= 22'h0101010001011100000010;
                12'h00d0: douta_buf <= 22'h1001010001011100000010;
                12'h00d1: douta_buf <= 22'h0001101001110100000010;
                12'h00d2: douta_buf <= 22'h0110000010001100000010;
                12'h00d3: douta_buf <= 22'h1010000010001100000010;
                12'h00d4: douta_buf <= 22'h0010011010100100000010;
                12'h00d5: douta_buf <= 22'h0110110010111100000010;
                12'h00d6: douta_buf <= 22'h1010110010111100000010;
                12'h00d7: douta_buf <= 22'h0000001000010100100110;
                12'h00d8: douta_buf <= 22'h0100100000101100100110;
                12'h00d9: douta_buf <= 22'h1000100000101100100110;
                12'h00da: douta_buf <= 22'h0000111001000100100110;
                12'h00db: douta_buf <= 22'h0101010001011100100110;
                12'h00dc: douta_buf <= 22'h1001010001011100100110;
                12'h00dd: douta_buf <= 22'h0001101001110100100110;
                12'h00de: douta_buf <= 22'h0110000010001100100110;
                12'h00df: douta_buf <= 22'h1010000010001100100110;
                12'h00e0: douta_buf <= 22'h0010011010100100100110;
                12'h00e1: douta_buf <= 22'h0110110010111100100110;
                12'h00e2: douta_buf <= 22'h1010110010111100100110;
                12'h00e3: douta_buf <= 22'h0001100000000000000001;
                12'h00e4: douta_buf <= 22'h0000000000000000000000;
                12'h00e5: douta_buf <= 22'h0000000000000000000000;
                12'h00e6: douta_buf <= 22'h0000000000000000000000;
                12'h00e7: douta_buf <= 22'h0000000000000000000000;
                12'h00e8: douta_buf <= 22'h0000000000001100000110;
                12'h00e9: douta_buf <= 22'h0000011000100100000110;
                12'h00ea: douta_buf <= 22'h0000110000111100000110;
                12'h00eb: douta_buf <= 22'h0001001001010100000110;
                12'h00ec: douta_buf <= 22'h0001100001101100000110;
                12'h00ed: douta_buf <= 22'h0001111010000100000110;
                12'h00ee: douta_buf <= 22'h0010010010011100000110;
                12'h00ef: douta_buf <= 22'h0010101010110100000110;
                12'h00f0: douta_buf <= 22'h0000000000001100100010;
                12'h00f1: douta_buf <= 22'h0000011000100100100010;
                12'h00f2: douta_buf <= 22'h0000110000111100100010;
                12'h00f3: douta_buf <= 22'h0001001001010100100010;
                12'h00f4: douta_buf <= 22'h0001100001101100100010;
                12'h00f5: douta_buf <= 22'h0001111010000100100010;
                12'h00f6: douta_buf <= 22'h0010010010011100100010;
                12'h00f7: douta_buf <= 22'h0010101010110100100010;
                12'h00f8: douta_buf <= 22'h0000000000001101001110;
                12'h00f9: douta_buf <= 22'h0000011000100101001110;
                12'h00fa: douta_buf <= 22'h0000110000111101001110;
                12'h00fb: douta_buf <= 22'h0001001001010101001110;
                12'h00fc: douta_buf <= 22'h0001100001101101001110;
                12'h00fd: douta_buf <= 22'h0001111010000101001110;
                12'h00fe: douta_buf <= 22'h0010010010011101001110;
                12'h00ff: douta_buf <= 22'h0010101010110101001110;
                12'h0100: douta_buf <= 22'h0000000000001101101010;
                12'h0101: douta_buf <= 22'h0000011000100101101010;
                12'h0102: douta_buf <= 22'h0000110000111101101010;
                12'h0103: douta_buf <= 22'h0001001001010101101010;
                12'h0104: douta_buf <= 22'h0001100001101101101010;
                12'h0105: douta_buf <= 22'h0001111010000101101010;
                12'h0106: douta_buf <= 22'h0010010010011101101010;
                12'h0107: douta_buf <= 22'h0010101010110101101010;
                12'h0108: douta_buf <= 22'h0000000100010000000110;
                12'h0109: douta_buf <= 22'h0000011100101000000110;
                12'h010a: douta_buf <= 22'h0000110101000000000110;
                12'h010b: douta_buf <= 22'h0001001101011000000110;
                12'h010c: douta_buf <= 22'h0001100101110000000110;
                12'h010d: douta_buf <= 22'h0001111110001000000110;
                12'h010e: douta_buf <= 22'h0010010110100000000110;
                12'h010f: douta_buf <= 22'h0010101110111000000110;
                12'h0110: douta_buf <= 22'h0000000100010000100010;
                12'h0111: douta_buf <= 22'h0000011100101000100010;
                12'h0112: douta_buf <= 22'h0000110101000000100010;
                12'h0113: douta_buf <= 22'h0001001101011000100010;
                12'h0114: douta_buf <= 22'h0001100101110000100010;
                12'h0115: douta_buf <= 22'h0001111110001000100010;
                12'h0116: douta_buf <= 22'h0010010110100000100010;
                12'h0117: douta_buf <= 22'h0010101110111000100010;
                12'h0118: douta_buf <= 22'h0000000100010001001110;
                12'h0119: douta_buf <= 22'h0000011100101001001110;
                12'h011a: douta_buf <= 22'h0000110101000001001110;
                12'h011b: douta_buf <= 22'h0001001101011001001110;
                12'h011c: douta_buf <= 22'h0001100101110001001110;
                12'h011d: douta_buf <= 22'h0001111110001001001110;
                12'h011e: douta_buf <= 22'h0010010110100001001110;
                12'h011f: douta_buf <= 22'h0010101110111001001110;
                12'h0120: douta_buf <= 22'h0000000100010001101010;
                12'h0121: douta_buf <= 22'h0000011100101001101010;
                12'h0122: douta_buf <= 22'h0000110101000001101010;
                12'h0123: douta_buf <= 22'h0001001101011001101010;
                12'h0124: douta_buf <= 22'h0001100101110001101010;
                12'h0125: douta_buf <= 22'h0001111110001001101010;
                12'h0126: douta_buf <= 22'h0010010110100001101010;
                12'h0127: douta_buf <= 22'h0010101110111001101010;
                12'h0128: douta_buf <= 22'h0000001000010100000110;
                12'h0129: douta_buf <= 22'h0000100000101100000110;
                12'h012a: douta_buf <= 22'h0000111001000100000110;
                12'h012b: douta_buf <= 22'h0001010001011100000110;
                12'h012c: douta_buf <= 22'h0001101001110100000110;
                12'h012d: douta_buf <= 22'h0010000010001100000110;
                12'h012e: douta_buf <= 22'h0010011010100100000110;
                12'h012f: douta_buf <= 22'h0010110010111100000110;
                12'h0130: douta_buf <= 22'h0000001000010100100010;
                12'h0131: douta_buf <= 22'h0000100000101100100010;
                12'h0132: douta_buf <= 22'h0000111001000100100010;
                12'h0133: douta_buf <= 22'h0001010001011100100010;
                12'h0134: douta_buf <= 22'h0001101001110100100010;
                12'h0135: douta_buf <= 22'h0010000010001100100010;
                12'h0136: douta_buf <= 22'h0010011010100100100010;
                12'h0137: douta_buf <= 22'h0010110010111100100010;
                12'h0138: douta_buf <= 22'h0000001000010101001110;
                12'h0139: douta_buf <= 22'h0000100000101101001110;
                12'h013a: douta_buf <= 22'h0000111001000101001110;
                12'h013b: douta_buf <= 22'h0001010001011101001110;
                12'h013c: douta_buf <= 22'h0001101001110101001110;
                12'h013d: douta_buf <= 22'h0010000010001101001110;
                12'h013e: douta_buf <= 22'h0010011010100101001110;
                12'h013f: douta_buf <= 22'h0010110010111101001110;
                12'h0140: douta_buf <= 22'h0000001000010101101010;
                12'h0141: douta_buf <= 22'h0000100000101101101010;
                12'h0142: douta_buf <= 22'h0000111001000101101010;
                12'h0143: douta_buf <= 22'h0001010001011101101010;
                12'h0144: douta_buf <= 22'h0001101001110101101010;
                12'h0145: douta_buf <= 22'h0010000010001101101010;
                12'h0146: douta_buf <= 22'h0010011010100101101010;
                12'h0147: douta_buf <= 22'h0010110010111101101010;
                12'h0148: douta_buf <= 22'h0001100000000000000001;
                12'h0149: douta_buf <= 22'h0000000000000000000000;
                12'h014a: douta_buf <= 22'h0000000000000000000000;
                12'h014b: douta_buf <= 22'h0000000000000000000000;
                12'h014c: douta_buf <= 22'h0000000000000000000000;
                12'h014d: douta_buf <= 22'h0000000000001100000110;
                12'h014e: douta_buf <= 22'h0100011000100100000110;
                12'h014f: douta_buf <= 22'h1000011000100100000110;
                12'h0150: douta_buf <= 22'h0000110000111100000110;
                12'h0151: douta_buf <= 22'h0101001001010100000110;
                12'h0152: douta_buf <= 22'h1001001001010100000110;
                12'h0153: douta_buf <= 22'h0001100001101100000110;
                12'h0154: douta_buf <= 22'h0101111010000100000110;
                12'h0155: douta_buf <= 22'h1001111010000100000110;
                12'h0156: douta_buf <= 22'h0010010010011100000110;
                12'h0157: douta_buf <= 22'h0110101010110100000110;
                12'h0158: douta_buf <= 22'h1010101010110100000110;
                12'h0159: douta_buf <= 22'h0000000000001100100010;
                12'h015a: douta_buf <= 22'h0100011000100100100010;
                12'h015b: douta_buf <= 22'h1000011000100100100010;
                12'h015c: douta_buf <= 22'h0000110000111100100010;
                12'h015d: douta_buf <= 22'h0101001001010100100010;
                12'h015e: douta_buf <= 22'h1001001001010100100010;
                12'h015f: douta_buf <= 22'h0001100001101100100010;
                12'h0160: douta_buf <= 22'h0101111010000100100010;
                12'h0161: douta_buf <= 22'h1001111010000100100010;
                12'h0162: douta_buf <= 22'h0010010010011100100010;
                12'h0163: douta_buf <= 22'h0110101010110100100010;
                12'h0164: douta_buf <= 22'h1010101010110100100010;
                12'h0165: douta_buf <= 22'h0000000000001101001110;
                12'h0166: douta_buf <= 22'h0100011000100101001110;
                12'h0167: douta_buf <= 22'h1000011000100101001110;
                12'h0168: douta_buf <= 22'h0000110000111101001110;
                12'h0169: douta_buf <= 22'h0101001001010101001110;
                12'h016a: douta_buf <= 22'h1001001001010101001110;
                12'h016b: douta_buf <= 22'h0001100001101101001110;
                12'h016c: douta_buf <= 22'h0101111010000101001110;
                12'h016d: douta_buf <= 22'h1001111010000101001110;
                12'h016e: douta_buf <= 22'h0010010010011101001110;
                12'h016f: douta_buf <= 22'h0110101010110101001110;
                12'h0170: douta_buf <= 22'h1010101010110101001110;
                12'h0171: douta_buf <= 22'h0000000000001101101010;
                12'h0172: douta_buf <= 22'h0100011000100101101010;
                12'h0173: douta_buf <= 22'h1000011000100101101010;
                12'h0174: douta_buf <= 22'h0000110000111101101010;
                12'h0175: douta_buf <= 22'h0101001001010101101010;
                12'h0176: douta_buf <= 22'h1001001001010101101010;
                12'h0177: douta_buf <= 22'h0001100001101101101010;
                12'h0178: douta_buf <= 22'h0101111010000101101010;
                12'h0179: douta_buf <= 22'h1001111010000101101010;
                12'h017a: douta_buf <= 22'h0010010010011101101010;
                12'h017b: douta_buf <= 22'h0110101010110101101010;
                12'h017c: douta_buf <= 22'h1010101010110101101010;
                12'h017d: douta_buf <= 22'h0000000100010000000110;
                12'h017e: douta_buf <= 22'h0100011100101000000110;
                12'h017f: douta_buf <= 22'h1000011100101000000110;
                12'h0180: douta_buf <= 22'h0000110101000000000110;
                12'h0181: douta_buf <= 22'h0101001101011000000110;
                12'h0182: douta_buf <= 22'h1001001101011000000110;
                12'h0183: douta_buf <= 22'h0001100101110000000110;
                12'h0184: douta_buf <= 22'h0101111110001000000110;
                12'h0185: douta_buf <= 22'h1001111110001000000110;
                12'h0186: douta_buf <= 22'h0010010110100000000110;
                12'h0187: douta_buf <= 22'h0110101110111000000110;
                12'h0188: douta_buf <= 22'h1010101110111000000110;
                12'h0189: douta_buf <= 22'h0000000100010000100010;
                12'h018a: douta_buf <= 22'h0100011100101000100010;
                12'h018b: douta_buf <= 22'h1000011100101000100010;
                12'h018c: douta_buf <= 22'h0000110101000000100010;
                12'h018d: douta_buf <= 22'h0101001101011000100010;
                12'h018e: douta_buf <= 22'h1001001101011000100010;
                12'h018f: douta_buf <= 22'h0001100101110000100010;
                12'h0190: douta_buf <= 22'h0101111110001000100010;
                12'h0191: douta_buf <= 22'h1001111110001000100010;
                12'h0192: douta_buf <= 22'h0010010110100000100010;
                12'h0193: douta_buf <= 22'h0110101110111000100010;
                12'h0194: douta_buf <= 22'h1010101110111000100010;
                12'h0195: douta_buf <= 22'h0000000100010001001110;
                12'h0196: douta_buf <= 22'h0100011100101001001110;
                12'h0197: douta_buf <= 22'h1000011100101001001110;
                12'h0198: douta_buf <= 22'h0000110101000001001110;
                12'h0199: douta_buf <= 22'h0101001101011001001110;
                12'h019a: douta_buf <= 22'h1001001101011001001110;
                12'h019b: douta_buf <= 22'h0001100101110001001110;
                12'h019c: douta_buf <= 22'h0101111110001001001110;
                12'h019d: douta_buf <= 22'h1001111110001001001110;
                12'h019e: douta_buf <= 22'h0010010110100001001110;
                12'h019f: douta_buf <= 22'h0110101110111001001110;
                12'h01a0: douta_buf <= 22'h1010101110111001001110;
                12'h01a1: douta_buf <= 22'h0000000100010001101010;
                12'h01a2: douta_buf <= 22'h0100011100101001101010;
                12'h01a3: douta_buf <= 22'h1000011100101001101010;
                12'h01a4: douta_buf <= 22'h0000110101000001101010;
                12'h01a5: douta_buf <= 22'h0101001101011001101010;
                12'h01a6: douta_buf <= 22'h1001001101011001101010;
                12'h01a7: douta_buf <= 22'h0001100101110001101010;
                12'h01a8: douta_buf <= 22'h0101111110001001101010;
                12'h01a9: douta_buf <= 22'h1001111110001001101010;
                12'h01aa: douta_buf <= 22'h0010010110100001101010;
                12'h01ab: douta_buf <= 22'h0110101110111001101010;
                12'h01ac: douta_buf <= 22'h1010101110111001101010;
                12'h01ad: douta_buf <= 22'h0000001000010100000110;
                12'h01ae: douta_buf <= 22'h0100100000101100000110;
                12'h01af: douta_buf <= 22'h1000100000101100000110;
                12'h01b0: douta_buf <= 22'h0000111001000100000110;
                12'h01b1: douta_buf <= 22'h0101010001011100000110;
                12'h01b2: douta_buf <= 22'h1001010001011100000110;
                12'h01b3: douta_buf <= 22'h0001101001110100000110;
                12'h01b4: douta_buf <= 22'h0110000010001100000110;
                12'h01b5: douta_buf <= 22'h1010000010001100000110;
                12'h01b6: douta_buf <= 22'h0010011010100100000110;
                12'h01b7: douta_buf <= 22'h0110110010111100000110;
                12'h01b8: douta_buf <= 22'h1010110010111100000110;
                12'h01b9: douta_buf <= 22'h0000001000010100100010;
                12'h01ba: douta_buf <= 22'h0100100000101100100010;
                12'h01bb: douta_buf <= 22'h1000100000101100100010;
                12'h01bc: douta_buf <= 22'h0000111001000100100010;
                12'h01bd: douta_buf <= 22'h0101010001011100100010;
                12'h01be: douta_buf <= 22'h1001010001011100100010;
                12'h01bf: douta_buf <= 22'h0001101001110100100010;
                12'h01c0: douta_buf <= 22'h0110000010001100100010;
                12'h01c1: douta_buf <= 22'h1010000010001100100010;
                12'h01c2: douta_buf <= 22'h0010011010100100100010;
                12'h01c3: douta_buf <= 22'h0110110010111100100010;
                12'h01c4: douta_buf <= 22'h1010110010111100100010;
                12'h01c5: douta_buf <= 22'h0000001000010101001110;
                12'h01c6: douta_buf <= 22'h0100100000101101001110;
                12'h01c7: douta_buf <= 22'h1000100000101101001110;
                12'h01c8: douta_buf <= 22'h0000111001000101001110;
                12'h01c9: douta_buf <= 22'h0101010001011101001110;
                12'h01ca: douta_buf <= 22'h1001010001011101001110;
                12'h01cb: douta_buf <= 22'h0001101001110101001110;
                12'h01cc: douta_buf <= 22'h0110000010001101001110;
                12'h01cd: douta_buf <= 22'h1010000010001101001110;
                12'h01ce: douta_buf <= 22'h0010011010100101001110;
                12'h01cf: douta_buf <= 22'h0110110010111101001110;
                12'h01d0: douta_buf <= 22'h1010110010111101001110;
                12'h01d1: douta_buf <= 22'h0000001000010101101010;
                12'h01d2: douta_buf <= 22'h0100100000101101101010;
                12'h01d3: douta_buf <= 22'h1000100000101101101010;
                12'h01d4: douta_buf <= 22'h0000111001000101101010;
                12'h01d5: douta_buf <= 22'h0101010001011101101010;
                12'h01d6: douta_buf <= 22'h1001010001011101101010;
                12'h01d7: douta_buf <= 22'h0001101001110101101010;
                12'h01d8: douta_buf <= 22'h0110000010001101101010;
                12'h01d9: douta_buf <= 22'h1010000010001101101010;
                12'h01da: douta_buf <= 22'h0010011010100101101010;
                12'h01db: douta_buf <= 22'h0110110010111101101010;
                12'h01dc: douta_buf <= 22'h1010110010111101101010;
                12'h01dd: douta_buf <= 22'h0001100000000000000001;
                12'h01de: douta_buf <= 22'h0000000000000000000000;
                12'h01df: douta_buf <= 22'h0000000000000000000000;
                12'h01e0: douta_buf <= 22'h0000000000000000000000;
                12'h01e1: douta_buf <= 22'h0000000000000000000000;
                12'h01e2: douta_buf <= 22'h0000000000001100001010;
                12'h01e3: douta_buf <= 22'h0100011000100100100010;
                12'h01e4: douta_buf <= 22'h0000100100110000001010;
                12'h01e5: douta_buf <= 22'h0100111101001000100010;
                12'h01e6: douta_buf <= 22'h0001001001010100001010;
                12'h01e7: douta_buf <= 22'h0101100001101100100010;
                12'h01e8: douta_buf <= 22'h0001101101111000001010;
                12'h01e9: douta_buf <= 22'h0110000110010000100010;
                12'h01ea: douta_buf <= 22'h0010010010011100001010;
                12'h01eb: douta_buf <= 22'h0110101010110100100010;
                12'h01ec: douta_buf <= 22'h0010110100000000000110;
                12'h01ed: douta_buf <= 22'h0100001100011000001010;
                12'h01ee: douta_buf <= 22'h0000011000100101000110;
                12'h01ef: douta_buf <= 22'h0100110000111100001010;
                12'h01f0: douta_buf <= 22'h0000111101001001000110;
                12'h01f1: douta_buf <= 22'h0101010101100000001010;
                12'h01f2: douta_buf <= 22'h0001100001101101000110;
                12'h01f3: douta_buf <= 22'h0101111010000100001010;
                12'h01f4: douta_buf <= 22'h0010000110010001000110;
                12'h01f5: douta_buf <= 22'h0110011110101000001010;
                12'h01f6: douta_buf <= 22'h0010101010110101000110;
                12'h01f7: douta_buf <= 22'h0100000000001101000110;
                12'h01f8: douta_buf <= 22'h0000001100011000100010;
                12'h01f9: douta_buf <= 22'h0100100100110001000110;
                12'h01fa: douta_buf <= 22'h0000110000111100100010;
                12'h01fb: douta_buf <= 22'h0101001001010101000110;
                12'h01fc: douta_buf <= 22'h0001010101100000100010;
                12'h01fd: douta_buf <= 22'h0101101101111001000110;
                12'h01fe: douta_buf <= 22'h0001111010000100100010;
                12'h01ff: douta_buf <= 22'h0110010010011101000110;
                12'h0200: douta_buf <= 22'h0010011110101000100010;
                12'h0201: douta_buf <= 22'h0110110100000001001110;
                12'h0202: douta_buf <= 22'h0000000000001101110110;
                12'h0203: douta_buf <= 22'h0100011000100110001110;
                12'h0204: douta_buf <= 22'h0000100100110001110110;
                12'h0205: douta_buf <= 22'h0100111101001010001110;
                12'h0206: douta_buf <= 22'h0001001001010101110110;
                12'h0207: douta_buf <= 22'h0101100001101110001110;
                12'h0208: douta_buf <= 22'h0001101101111001110110;
                12'h0209: douta_buf <= 22'h0110000110010010001110;
                12'h020a: douta_buf <= 22'h0010010010011101110110;
                12'h020b: douta_buf <= 22'h0110101010110110001110;
                12'h020c: douta_buf <= 22'h0010110100000001110010;
                12'h020d: douta_buf <= 22'h0100001100011001110110;
                12'h020e: douta_buf <= 22'h0000011000100110110010;
                12'h020f: douta_buf <= 22'h0100110000111101110110;
                12'h0210: douta_buf <= 22'h0000111101001010110010;
                12'h0211: douta_buf <= 22'h0101010101100001110110;
                12'h0212: douta_buf <= 22'h0001100001101110110010;
                12'h0213: douta_buf <= 22'h0101111010000101110110;
                12'h0214: douta_buf <= 22'h0010000110010010110010;
                12'h0215: douta_buf <= 22'h0110011110101001110110;
                12'h0216: douta_buf <= 22'h0010101010110110110010;
                12'h0217: douta_buf <= 22'h0100000000001110110010;
                12'h0218: douta_buf <= 22'h0000001100011010001110;
                12'h0219: douta_buf <= 22'h0100100100110010110010;
                12'h021a: douta_buf <= 22'h0000110000111110001110;
                12'h021b: douta_buf <= 22'h0101001001010110110010;
                12'h021c: douta_buf <= 22'h0001010101100010001110;
                12'h021d: douta_buf <= 22'h0101101101111010110010;
                12'h021e: douta_buf <= 22'h0001111010000110001110;
                12'h021f: douta_buf <= 22'h0110010010011110110010;
                12'h0220: douta_buf <= 22'h0010011110101010001110;
                12'h0221: douta_buf <= 22'h0110110100000110100010;
                12'h0222: douta_buf <= 22'h0000000100010000001010;
                12'h0223: douta_buf <= 22'h0100011100101000100010;
                12'h0224: douta_buf <= 22'h0000101000110100001010;
                12'h0225: douta_buf <= 22'h0101000001001100100010;
                12'h0226: douta_buf <= 22'h0001001101011000001010;
                12'h0227: douta_buf <= 22'h0101100101110000100010;
                12'h0228: douta_buf <= 22'h0001110001111100001010;
                12'h0229: douta_buf <= 22'h0110001010010100100010;
                12'h022a: douta_buf <= 22'h0010010110100000001010;
                12'h022b: douta_buf <= 22'h0110101110111000100010;
                12'h022c: douta_buf <= 22'h0010111000000100000110;
                12'h022d: douta_buf <= 22'h0100010000011100001010;
                12'h022e: douta_buf <= 22'h0000011100101001000110;
                12'h022f: douta_buf <= 22'h0100110101000000001010;
                12'h0230: douta_buf <= 22'h0001000001001101000110;
                12'h0231: douta_buf <= 22'h0101011001100100001010;
                12'h0232: douta_buf <= 22'h0001100101110001000110;
                12'h0233: douta_buf <= 22'h0101111110001000001010;
                12'h0234: douta_buf <= 22'h0010001010010101000110;
                12'h0235: douta_buf <= 22'h0110100010101100001010;
                12'h0236: douta_buf <= 22'h0010101110111001000110;
                12'h0237: douta_buf <= 22'h0100000100010001000110;
                12'h0238: douta_buf <= 22'h0000010000011100100010;
                12'h0239: douta_buf <= 22'h0100101000110101000110;
                12'h023a: douta_buf <= 22'h0000110101000000100010;
                12'h023b: douta_buf <= 22'h0101001101011001000110;
                12'h023c: douta_buf <= 22'h0001011001100100100010;
                12'h023d: douta_buf <= 22'h0101110001111101000110;
                12'h023e: douta_buf <= 22'h0001111110001000100010;
                12'h023f: douta_buf <= 22'h0110010110100001000110;
                12'h0240: douta_buf <= 22'h0010100010101100100010;
                12'h0241: douta_buf <= 22'h0110111000000101001110;
                12'h0242: douta_buf <= 22'h0000000100010001110110;
                12'h0243: douta_buf <= 22'h0100011100101010001110;
                12'h0244: douta_buf <= 22'h0000101000110101110110;
                12'h0245: douta_buf <= 22'h0101000001001110001110;
                12'h0246: douta_buf <= 22'h0001001101011001110110;
                12'h0247: douta_buf <= 22'h0101100101110010001110;
                12'h0248: douta_buf <= 22'h0001110001111101110110;
                12'h0249: douta_buf <= 22'h0110001010010110001110;
                12'h024a: douta_buf <= 22'h0010010110100001110110;
                12'h024b: douta_buf <= 22'h0110101110111010001110;
                12'h024c: douta_buf <= 22'h0010111000000101110010;
                12'h024d: douta_buf <= 22'h0100010000011101110110;
                12'h024e: douta_buf <= 22'h0000011100101010110010;
                12'h024f: douta_buf <= 22'h0100110101000001110110;
                12'h0250: douta_buf <= 22'h0001000001001110110010;
                12'h0251: douta_buf <= 22'h0101011001100101110110;
                12'h0252: douta_buf <= 22'h0001100101110010110010;
                12'h0253: douta_buf <= 22'h0101111110001001110110;
                12'h0254: douta_buf <= 22'h0010001010010110110010;
                12'h0255: douta_buf <= 22'h0110100010101101110110;
                12'h0256: douta_buf <= 22'h0010101110111010110010;
                12'h0257: douta_buf <= 22'h0100000100010010110010;
                12'h0258: douta_buf <= 22'h0000010000011110001110;
                12'h0259: douta_buf <= 22'h0100101000110110110010;
                12'h025a: douta_buf <= 22'h0000110101000010001110;
                12'h025b: douta_buf <= 22'h0101001101011010110010;
                12'h025c: douta_buf <= 22'h0001011001100110001110;
                12'h025d: douta_buf <= 22'h0101110001111110110010;
                12'h025e: douta_buf <= 22'h0001111110001010001110;
                12'h025f: douta_buf <= 22'h0110010110100010110010;
                12'h0260: douta_buf <= 22'h0010100010101110001110;
                12'h0261: douta_buf <= 22'h0110111000001010100010;
                12'h0262: douta_buf <= 22'h0000001000010100001010;
                12'h0263: douta_buf <= 22'h0100100000101100100010;
                12'h0264: douta_buf <= 22'h0000101100111000001010;
                12'h0265: douta_buf <= 22'h0101000101010000100010;
                12'h0266: douta_buf <= 22'h0001010001011100001010;
                12'h0267: douta_buf <= 22'h0101101001110100100010;
                12'h0268: douta_buf <= 22'h0001110110000000001010;
                12'h0269: douta_buf <= 22'h0110001110011000100010;
                12'h026a: douta_buf <= 22'h0010011010100100001010;
                12'h026b: douta_buf <= 22'h0110110010111100100010;
                12'h026c: douta_buf <= 22'h0010111100001000000110;
                12'h026d: douta_buf <= 22'h0100010100100000001010;
                12'h026e: douta_buf <= 22'h0000100000101101000110;
                12'h026f: douta_buf <= 22'h0100111001000100001010;
                12'h0270: douta_buf <= 22'h0001000101010001000110;
                12'h0271: douta_buf <= 22'h0101011101101000001010;
                12'h0272: douta_buf <= 22'h0001101001110101000110;
                12'h0273: douta_buf <= 22'h0110000010001100001010;
                12'h0274: douta_buf <= 22'h0010001110011001000110;
                12'h0275: douta_buf <= 22'h0110100110110000001010;
                12'h0276: douta_buf <= 22'h0010110010111101000110;
                12'h0277: douta_buf <= 22'h0100001000010101000110;
                12'h0278: douta_buf <= 22'h0000010100100000100010;
                12'h0279: douta_buf <= 22'h0100101100111001000110;
                12'h027a: douta_buf <= 22'h0000111001000100100010;
                12'h027b: douta_buf <= 22'h0101010001011101000110;
                12'h027c: douta_buf <= 22'h0001011101101000100010;
                12'h027d: douta_buf <= 22'h0101110110000001000110;
                12'h027e: douta_buf <= 22'h0010000010001100100010;
                12'h027f: douta_buf <= 22'h0110011010100101000110;
                12'h0280: douta_buf <= 22'h0010100110110000100010;
                12'h0281: douta_buf <= 22'h0110111100001001001110;
                12'h0282: douta_buf <= 22'h0000001000010101110110;
                12'h0283: douta_buf <= 22'h0100100000101110001110;
                12'h0284: douta_buf <= 22'h0000101100111001110110;
                12'h0285: douta_buf <= 22'h0101000101010010001110;
                12'h0286: douta_buf <= 22'h0001010001011101110110;
                12'h0287: douta_buf <= 22'h0101101001110110001110;
                12'h0288: douta_buf <= 22'h0001110110000001110110;
                12'h0289: douta_buf <= 22'h0110001110011010001110;
                12'h028a: douta_buf <= 22'h0010011010100101110110;
                12'h028b: douta_buf <= 22'h0110110010111110001110;
                12'h028c: douta_buf <= 22'h0010111100001001110010;
                12'h028d: douta_buf <= 22'h0100010100100001110110;
                12'h028e: douta_buf <= 22'h0000100000101110110010;
                12'h028f: douta_buf <= 22'h0100111001000101110110;
                12'h0290: douta_buf <= 22'h0001000101010010110010;
                12'h0291: douta_buf <= 22'h0101011101101001110110;
                12'h0292: douta_buf <= 22'h0001101001110110110010;
                12'h0293: douta_buf <= 22'h0110000010001101110110;
                12'h0294: douta_buf <= 22'h0010001110011010110010;
                12'h0295: douta_buf <= 22'h0110100110110001110110;
                12'h0296: douta_buf <= 22'h0010110010111110110010;
                12'h0297: douta_buf <= 22'h0100001000010110110010;
                12'h0298: douta_buf <= 22'h0000010100100010001110;
                12'h0299: douta_buf <= 22'h0100101100111010110010;
                12'h029a: douta_buf <= 22'h0000111001000110001110;
                12'h029b: douta_buf <= 22'h0101010001011110110010;
                12'h029c: douta_buf <= 22'h0001011101101010001110;
                12'h029d: douta_buf <= 22'h0101110110000010110010;
                12'h029e: douta_buf <= 22'h0010000010001110001110;
                12'h029f: douta_buf <= 22'h0110011010100110110010;
                12'h02a0: douta_buf <= 22'h0010100110110010001110;
                12'h02a1: douta_buf <= 22'h0110111100000010100010;
                12'h02a2: douta_buf <= 22'h0001100000000000000001;
                12'h02a3: douta_buf <= 22'h0000000000000000000000;
                12'h02a4: douta_buf <= 22'h0000000000000000000000;
                12'h02a5: douta_buf <= 22'h0000000000000000000000;
                12'h02a6: douta_buf <= 22'h0000000000000000000000;
                12'h02a7: douta_buf <= 22'h0000000000001100001010;
                12'h02a8: douta_buf <= 22'h0100011000100100100010;
                12'h02a9: douta_buf <= 22'h1000011000100100100010;
                12'h02aa: douta_buf <= 22'h0000110000111101000110;
                12'h02ab: douta_buf <= 22'h0101001001010100001010;
                12'h02ac: douta_buf <= 22'h1001001001010100001010;
                12'h02ad: douta_buf <= 22'h0001100001101100100010;
                12'h02ae: douta_buf <= 22'h0101111010000101000110;
                12'h02af: douta_buf <= 22'h1001111010000101000110;
                12'h02b0: douta_buf <= 22'h0010010010011100001010;
                12'h02b1: douta_buf <= 22'h0110101010110100100010;
                12'h02b2: douta_buf <= 22'h1010101010110100100010;
                12'h02b3: douta_buf <= 22'h0000000000001100100010;
                12'h02b4: douta_buf <= 22'h0100011000100101000110;
                12'h02b5: douta_buf <= 22'h1000011000100101000110;
                12'h02b6: douta_buf <= 22'h0000110000111100001010;
                12'h02b7: douta_buf <= 22'h0101001001010100100010;
                12'h02b8: douta_buf <= 22'h1001001001010100100010;
                12'h02b9: douta_buf <= 22'h0001100001101101000110;
                12'h02ba: douta_buf <= 22'h0101111010000100001010;
                12'h02bb: douta_buf <= 22'h1001111010000100001010;
                12'h02bc: douta_buf <= 22'h0010010010011100100010;
                12'h02bd: douta_buf <= 22'h0110101010110101000110;
                12'h02be: douta_buf <= 22'h1010101010110101000110;
                12'h02bf: douta_buf <= 22'h0000000000001101000110;
                12'h02c0: douta_buf <= 22'h0100011000100100001010;
                12'h02c1: douta_buf <= 22'h1000011000100100001010;
                12'h02c2: douta_buf <= 22'h0000110000111100100010;
                12'h02c3: douta_buf <= 22'h0101001001010101000110;
                12'h02c4: douta_buf <= 22'h1001001001010101000110;
                12'h02c5: douta_buf <= 22'h0001100001101100001010;
                12'h02c6: douta_buf <= 22'h0101111010000100100010;
                12'h02c7: douta_buf <= 22'h1001111010000100100010;
                12'h02c8: douta_buf <= 22'h0010010010011101000110;
                12'h02c9: douta_buf <= 22'h0110101010110100001010;
                12'h02ca: douta_buf <= 22'h1010101010110100001010;
                12'h02cb: douta_buf <= 22'h0000000000001101110110;
                12'h02cc: douta_buf <= 22'h0100011000100110001110;
                12'h02cd: douta_buf <= 22'h1000011000100110001110;
                12'h02ce: douta_buf <= 22'h0000110000111110110010;
                12'h02cf: douta_buf <= 22'h0101001001010101110110;
                12'h02d0: douta_buf <= 22'h1001001001010101110110;
                12'h02d1: douta_buf <= 22'h0001100001101110001110;
                12'h02d2: douta_buf <= 22'h0101111010000110110010;
                12'h02d3: douta_buf <= 22'h1001111010000110110010;
                12'h02d4: douta_buf <= 22'h0010010010011101110110;
                12'h02d5: douta_buf <= 22'h0110101010110110001110;
                12'h02d6: douta_buf <= 22'h1010101010110110001110;
                12'h02d7: douta_buf <= 22'h0000000000001110001110;
                12'h02d8: douta_buf <= 22'h0100011000100110110010;
                12'h02d9: douta_buf <= 22'h1000011000100110110010;
                12'h02da: douta_buf <= 22'h0000110000111101110110;
                12'h02db: douta_buf <= 22'h0101001001010110001110;
                12'h02dc: douta_buf <= 22'h1001001001010110001110;
                12'h02dd: douta_buf <= 22'h0001100001101110110010;
                12'h02de: douta_buf <= 22'h0101111010000101110110;
                12'h02df: douta_buf <= 22'h1001111010000101110110;
                12'h02e0: douta_buf <= 22'h0010010010011110001110;
                12'h02e1: douta_buf <= 22'h0110101010110110110010;
                12'h02e2: douta_buf <= 22'h1010101010110110110010;
                12'h02e3: douta_buf <= 22'h0000000000001110110010;
                12'h02e4: douta_buf <= 22'h0100011000100101110110;
                12'h02e5: douta_buf <= 22'h1000011000100101110110;
                12'h02e6: douta_buf <= 22'h0000110000111110001110;
                12'h02e7: douta_buf <= 22'h0101001001010110110010;
                12'h02e8: douta_buf <= 22'h1001001001010110110010;
                12'h02e9: douta_buf <= 22'h0001100001101101110110;
                12'h02ea: douta_buf <= 22'h0101111010000110001110;
                12'h02eb: douta_buf <= 22'h1001111010000110001110;
                12'h02ec: douta_buf <= 22'h0010010010011110110010;
                12'h02ed: douta_buf <= 22'h0110101010110101110110;
                12'h02ee: douta_buf <= 22'h1010101010110101110110;
                12'h02ef: douta_buf <= 22'h0000000100010000001010;
                12'h02f0: douta_buf <= 22'h0100011100101000100010;
                12'h02f1: douta_buf <= 22'h1000011100101000100010;
                12'h02f2: douta_buf <= 22'h0000110101000001000110;
                12'h02f3: douta_buf <= 22'h0101001101011000001010;
                12'h02f4: douta_buf <= 22'h1001001101011000001010;
                12'h02f5: douta_buf <= 22'h0001100101110000100010;
                12'h02f6: douta_buf <= 22'h0101111110001001000110;
                12'h02f7: douta_buf <= 22'h1001111110001001000110;
                12'h02f8: douta_buf <= 22'h0010010110100000001010;
                12'h02f9: douta_buf <= 22'h0110101110111000100010;
                12'h02fa: douta_buf <= 22'h1010101110111000100010;
                12'h02fb: douta_buf <= 22'h0000000100010000100010;
                12'h02fc: douta_buf <= 22'h0100011100101001000110;
                12'h02fd: douta_buf <= 22'h1000011100101001000110;
                12'h02fe: douta_buf <= 22'h0000110101000000001010;
                12'h02ff: douta_buf <= 22'h0101001101011000100010;
                12'h0300: douta_buf <= 22'h1001001101011000100010;
                12'h0301: douta_buf <= 22'h0001100101110001000110;
                12'h0302: douta_buf <= 22'h0101111110001000001010;
                12'h0303: douta_buf <= 22'h1001111110001000001010;
                12'h0304: douta_buf <= 22'h0010010110100000100010;
                12'h0305: douta_buf <= 22'h0110101110111001000110;
                12'h0306: douta_buf <= 22'h1010101110111001000110;
                12'h0307: douta_buf <= 22'h0000000100010001000110;
                12'h0308: douta_buf <= 22'h0100011100101000001010;
                12'h0309: douta_buf <= 22'h1000011100101000001010;
                12'h030a: douta_buf <= 22'h0000110101000000100010;
                12'h030b: douta_buf <= 22'h0101001101011001000110;
                12'h030c: douta_buf <= 22'h1001001101011001000110;
                12'h030d: douta_buf <= 22'h0001100101110000001010;
                12'h030e: douta_buf <= 22'h0101111110001000100010;
                12'h030f: douta_buf <= 22'h1001111110001000100010;
                12'h0310: douta_buf <= 22'h0010010110100001000110;
                12'h0311: douta_buf <= 22'h0110101110111000001010;
                12'h0312: douta_buf <= 22'h1010101110111000001010;
                12'h0313: douta_buf <= 22'h0000000100010001110110;
                12'h0314: douta_buf <= 22'h0100011100101010001110;
                12'h0315: douta_buf <= 22'h1000011100101010001110;
                12'h0316: douta_buf <= 22'h0000110101000010110010;
                12'h0317: douta_buf <= 22'h0101001101011001110110;
                12'h0318: douta_buf <= 22'h1001001101011001110110;
                12'h0319: douta_buf <= 22'h0001100101110010001110;
                12'h031a: douta_buf <= 22'h0101111110001010110010;
                12'h031b: douta_buf <= 22'h1001111110001010110010;
                12'h031c: douta_buf <= 22'h0010010110100001110110;
                12'h031d: douta_buf <= 22'h0110101110111010001110;
                12'h031e: douta_buf <= 22'h1010101110111010001110;
                12'h031f: douta_buf <= 22'h0000000100010010001110;
                12'h0320: douta_buf <= 22'h0100011100101010110010;
                12'h0321: douta_buf <= 22'h1000011100101010110010;
                12'h0322: douta_buf <= 22'h0000110101000001110110;
                12'h0323: douta_buf <= 22'h0101001101011010001110;
                12'h0324: douta_buf <= 22'h1001001101011010001110;
                12'h0325: douta_buf <= 22'h0001100101110010110010;
                12'h0326: douta_buf <= 22'h0101111110001001110110;
                12'h0327: douta_buf <= 22'h1001111110001001110110;
                12'h0328: douta_buf <= 22'h0010010110100010001110;
                12'h0329: douta_buf <= 22'h0110101110111010110010;
                12'h032a: douta_buf <= 22'h1010101110111010110010;
                12'h032b: douta_buf <= 22'h0000000100010010110010;
                12'h032c: douta_buf <= 22'h0100011100101001110110;
                12'h032d: douta_buf <= 22'h1000011100101001110110;
                12'h032e: douta_buf <= 22'h0000110101000010001110;
                12'h032f: douta_buf <= 22'h0101001101011010110010;
                12'h0330: douta_buf <= 22'h1001001101011010110010;
                12'h0331: douta_buf <= 22'h0001100101110001110110;
                12'h0332: douta_buf <= 22'h0101111110001010001110;
                12'h0333: douta_buf <= 22'h1001111110001010001110;
                12'h0334: douta_buf <= 22'h0010010110100010110010;
                12'h0335: douta_buf <= 22'h0110101110111001110110;
                12'h0336: douta_buf <= 22'h1010101110111001110110;
                12'h0337: douta_buf <= 22'h0000001000010100001010;
                12'h0338: douta_buf <= 22'h0100100000101100100010;
                12'h0339: douta_buf <= 22'h1000100000101100100010;
                12'h033a: douta_buf <= 22'h0000111001000101000110;
                12'h033b: douta_buf <= 22'h0101010001011100001010;
                12'h033c: douta_buf <= 22'h1001010001011100001010;
                12'h033d: douta_buf <= 22'h0001101001110100100010;
                12'h033e: douta_buf <= 22'h0110000010001101000110;
                12'h033f: douta_buf <= 22'h1010000010001101000110;
                12'h0340: douta_buf <= 22'h0010011010100100001010;
                12'h0341: douta_buf <= 22'h0110110010111100100010;
                12'h0342: douta_buf <= 22'h1010110010111100100010;
                12'h0343: douta_buf <= 22'h0000001000010100100010;
                12'h0344: douta_buf <= 22'h0100100000101101000110;
                12'h0345: douta_buf <= 22'h1000100000101101000110;
                12'h0346: douta_buf <= 22'h0000111001000100001010;
                12'h0347: douta_buf <= 22'h0101010001011100100010;
                12'h0348: douta_buf <= 22'h1001010001011100100010;
                12'h0349: douta_buf <= 22'h0001101001110101000110;
                12'h034a: douta_buf <= 22'h0110000010001100001010;
                12'h034b: douta_buf <= 22'h1010000010001100001010;
                12'h034c: douta_buf <= 22'h0010011010100100100010;
                12'h034d: douta_buf <= 22'h0110110010111101000110;
                12'h034e: douta_buf <= 22'h1010110010111101000110;
                12'h034f: douta_buf <= 22'h0000001000010101000110;
                12'h0350: douta_buf <= 22'h0100100000101100001010;
                12'h0351: douta_buf <= 22'h1000100000101100001010;
                12'h0352: douta_buf <= 22'h0000111001000100100010;
                12'h0353: douta_buf <= 22'h0101010001011101000110;
                12'h0354: douta_buf <= 22'h1001010001011101000110;
                12'h0355: douta_buf <= 22'h0001101001110100001010;
                12'h0356: douta_buf <= 22'h0110000010001100100010;
                12'h0357: douta_buf <= 22'h1010000010001100100010;
                12'h0358: douta_buf <= 22'h0010011010100101000110;
                12'h0359: douta_buf <= 22'h0110110010111100001010;
                12'h035a: douta_buf <= 22'h1010110010111100001010;
                12'h035b: douta_buf <= 22'h0000001000010101110110;
                12'h035c: douta_buf <= 22'h0100100000101110001110;
                12'h035d: douta_buf <= 22'h1000100000101110001110;
                12'h035e: douta_buf <= 22'h0000111001000110110010;
                12'h035f: douta_buf <= 22'h0101010001011101110110;
                12'h0360: douta_buf <= 22'h1001010001011101110110;
                12'h0361: douta_buf <= 22'h0001101001110110001110;
                12'h0362: douta_buf <= 22'h0110000010001110110010;
                12'h0363: douta_buf <= 22'h1010000010001110110010;
                12'h0364: douta_buf <= 22'h0010011010100101110110;
                12'h0365: douta_buf <= 22'h0110110010111110001110;
                12'h0366: douta_buf <= 22'h1010110010111110001110;
                12'h0367: douta_buf <= 22'h0000001000010110001110;
                12'h0368: douta_buf <= 22'h0100100000101110110010;
                12'h0369: douta_buf <= 22'h1000100000101110110010;
                12'h036a: douta_buf <= 22'h0000111001000101110110;
                12'h036b: douta_buf <= 22'h0101010001011110001110;
                12'h036c: douta_buf <= 22'h1001010001011110001110;
                12'h036d: douta_buf <= 22'h0001101001110110110010;
                12'h036e: douta_buf <= 22'h0110000010001101110110;
                12'h036f: douta_buf <= 22'h1010000010001101110110;
                12'h0370: douta_buf <= 22'h0010011010100110001110;
                12'h0371: douta_buf <= 22'h0110110010111110110010;
                12'h0372: douta_buf <= 22'h1010110010111110110010;
                12'h0373: douta_buf <= 22'h0000001000010110110010;
                12'h0374: douta_buf <= 22'h0100100000101101110110;
                12'h0375: douta_buf <= 22'h1000100000101101110110;
                12'h0376: douta_buf <= 22'h0000111001000110001110;
                12'h0377: douta_buf <= 22'h0101010001011110110010;
                12'h0378: douta_buf <= 22'h1001010001011110110010;
                12'h0379: douta_buf <= 22'h0001101001110101110110;
                12'h037a: douta_buf <= 22'h0110000010001110001110;
                12'h037b: douta_buf <= 22'h1010000010001110001110;
                12'h037c: douta_buf <= 22'h0010011010100110110010;
                12'h037d: douta_buf <= 22'h0110110010111101110110;
                12'h037e: douta_buf <= 22'h1010110010111101110110;
                12'h037f: douta_buf <= 22'h0001100000000000000001;
                12'h0380: douta_buf <= 22'h0000000000000000000000;
                12'h0381: douta_buf <= 22'h0000000000000000000000;
                12'h0382: douta_buf <= 22'h0000000000000000000000;
                12'h0383: douta_buf <= 22'h0000000000000000000000;
                12'h0384: douta_buf <= 22'h0000000000010000000010;
                12'h0385: douta_buf <= 22'h0000100000110000000010;
                12'h0386: douta_buf <= 22'h0001000001010000000010;
                12'h0387: douta_buf <= 22'h0001100001110000000010;
                12'h0388: douta_buf <= 22'h0010000010010000000010;
                12'h0389: douta_buf <= 22'h0010100010110000000010;
                12'h038a: douta_buf <= 22'h0011000000000100000010;
                12'h038b: douta_buf <= 22'h0000010100100100000010;
                12'h038c: douta_buf <= 22'h0000110101000100000010;
                12'h038d: douta_buf <= 22'h0001010101100100000010;
                12'h038e: douta_buf <= 22'h0001110110000100000010;
                12'h038f: douta_buf <= 22'h0010010110100100000010;
                12'h0390: douta_buf <= 22'h0010110111000100000010;
                12'h0391: douta_buf <= 22'h0000001000011000000010;
                12'h0392: douta_buf <= 22'h0000101000111000000010;
                12'h0393: douta_buf <= 22'h0001001001011000000010;
                12'h0394: douta_buf <= 22'h0001101001111000000010;
                12'h0395: douta_buf <= 22'h0010001010011000000010;
                12'h0396: douta_buf <= 22'h0010101010111000000010;
                12'h0397: douta_buf <= 22'h0011001000001100000010;
                12'h0398: douta_buf <= 22'h0000011100101100000010;
                12'h0399: douta_buf <= 22'h0000111101001100000010;
                12'h039a: douta_buf <= 22'h0001011101101100000010;
                12'h039b: douta_buf <= 22'h0001111110001100000010;
                12'h039c: douta_buf <= 22'h0010011110101100000010;
                12'h039d: douta_buf <= 22'h0010111111001100000010;
                12'h039e: douta_buf <= 22'h0001101000000000000001;
                12'h039f: douta_buf <= 22'h0000000000000000000000;
                12'h03a0: douta_buf <= 22'h0000000000000000000000;
                12'h03a1: douta_buf <= 22'h0000000000000000000000;
                12'h03a2: douta_buf <= 22'h0000000000000000000000;
                12'h03a3: douta_buf <= 22'h0000000000010000000010;
                12'h03a4: douta_buf <= 22'h0000100000110000000010;
                12'h03a5: douta_buf <= 22'h0001000001010000000010;
                12'h03a6: douta_buf <= 22'h0001100001110000000010;
                12'h03a7: douta_buf <= 22'h0010000010010000000010;
                12'h03a8: douta_buf <= 22'h0010100010110000000010;
                12'h03a9: douta_buf <= 22'h0011000000000000000110;
                12'h03aa: douta_buf <= 22'h0000010000100000100110;
                12'h03ab: douta_buf <= 22'h0000110001000000100110;
                12'h03ac: douta_buf <= 22'h0001010001100000100110;
                12'h03ad: douta_buf <= 22'h0001110010000000100110;
                12'h03ae: douta_buf <= 22'h0010010010100000100110;
                12'h03af: douta_buf <= 22'h0010110011000000100110;
                12'h03b0: douta_buf <= 22'h0000000100010100000010;
                12'h03b1: douta_buf <= 22'h0000100100110100000010;
                12'h03b2: douta_buf <= 22'h0001000101010100000010;
                12'h03b3: douta_buf <= 22'h0001100101110100000010;
                12'h03b4: douta_buf <= 22'h0010000110010100000010;
                12'h03b5: douta_buf <= 22'h0010100110110100000010;
                12'h03b6: douta_buf <= 22'h0011000100000100000110;
                12'h03b7: douta_buf <= 22'h0000010100100100100110;
                12'h03b8: douta_buf <= 22'h0000110101000100100110;
                12'h03b9: douta_buf <= 22'h0001010101100100100110;
                12'h03ba: douta_buf <= 22'h0001110110000100100110;
                12'h03bb: douta_buf <= 22'h0010010110100100100110;
                12'h03bc: douta_buf <= 22'h0010110111000100100110;
                12'h03bd: douta_buf <= 22'h0000001000011000000010;
                12'h03be: douta_buf <= 22'h0000101000111000000010;
                12'h03bf: douta_buf <= 22'h0001001001011000000010;
                12'h03c0: douta_buf <= 22'h0001101001111000000010;
                12'h03c1: douta_buf <= 22'h0010001010011000000010;
                12'h03c2: douta_buf <= 22'h0010101010111000000010;
                12'h03c3: douta_buf <= 22'h0011001000001000000110;
                12'h03c4: douta_buf <= 22'h0000011000101000100110;
                12'h03c5: douta_buf <= 22'h0000111001001000100110;
                12'h03c6: douta_buf <= 22'h0001011001101000100110;
                12'h03c7: douta_buf <= 22'h0001111010001000100110;
                12'h03c8: douta_buf <= 22'h0010011010101000100110;
                12'h03c9: douta_buf <= 22'h0010111011001000100110;
                12'h03ca: douta_buf <= 22'h0000001100011100000010;
                12'h03cb: douta_buf <= 22'h0000101100111100000010;
                12'h03cc: douta_buf <= 22'h0001001101011100000010;
                12'h03cd: douta_buf <= 22'h0001101101111100000010;
                12'h03ce: douta_buf <= 22'h0010001110011100000010;
                12'h03cf: douta_buf <= 22'h0010101110111100000010;
                12'h03d0: douta_buf <= 22'h0011001100001100000110;
                12'h03d1: douta_buf <= 22'h0000011100101100100110;
                12'h03d2: douta_buf <= 22'h0000111101001100100110;
                12'h03d3: douta_buf <= 22'h0001011101101100100110;
                12'h03d4: douta_buf <= 22'h0001111110001100100110;
                12'h03d5: douta_buf <= 22'h0010011110101100100110;
                12'h03d6: douta_buf <= 22'h0010111111001100100110;
                12'h03d7: douta_buf <= 22'h0001101000000000000001;
                12'h03d8: douta_buf <= 22'h0000000000000000000000;
                12'h03d9: douta_buf <= 22'h0000000000000000000000;
                12'h03da: douta_buf <= 22'h0000000000000000000000;
                12'h03db: douta_buf <= 22'h0000000000000000000000;
                12'h03dc: douta_buf <= 22'h0000000000010000000010;
                12'h03dd: douta_buf <= 22'h0100100000110000000010;
                12'h03de: douta_buf <= 22'h1000100000110000000010;
                12'h03df: douta_buf <= 22'h0001000001010000000010;
                12'h03e0: douta_buf <= 22'h0101100001110000000010;
                12'h03e1: douta_buf <= 22'h1001100001110000000010;
                12'h03e2: douta_buf <= 22'h0010000010010000000010;
                12'h03e3: douta_buf <= 22'h0110100010110000000010;
                12'h03e4: douta_buf <= 22'h1010100010110000000010;
                12'h03e5: douta_buf <= 22'h0011000000000000000110;
                12'h03e6: douta_buf <= 22'h0100010000100000100110;
                12'h03e7: douta_buf <= 22'h1000010000100000100110;
                12'h03e8: douta_buf <= 22'h0000110001000000100110;
                12'h03e9: douta_buf <= 22'h0101010001100000100110;
                12'h03ea: douta_buf <= 22'h1001010001100000100110;
                12'h03eb: douta_buf <= 22'h0001110010000000100110;
                12'h03ec: douta_buf <= 22'h0110010010100000100110;
                12'h03ed: douta_buf <= 22'h1010010010100000100110;
                12'h03ee: douta_buf <= 22'h0010110011000000100110;
                12'h03ef: douta_buf <= 22'h0100000100010100000010;
                12'h03f0: douta_buf <= 22'h1000000100010100000010;
                12'h03f1: douta_buf <= 22'h0000100100110100000010;
                12'h03f2: douta_buf <= 22'h0101000101010100000010;
                12'h03f3: douta_buf <= 22'h1001000101010100000010;
                12'h03f4: douta_buf <= 22'h0001100101110100000010;
                12'h03f5: douta_buf <= 22'h0110000110010100000010;
                12'h03f6: douta_buf <= 22'h1010000110010100000010;
                12'h03f7: douta_buf <= 22'h0010100110110100000010;
                12'h03f8: douta_buf <= 22'h0111000100000100000110;
                12'h03f9: douta_buf <= 22'h1011000100000100000110;
                12'h03fa: douta_buf <= 22'h0000010100100100100110;
                12'h03fb: douta_buf <= 22'h0100110101000100100110;
                12'h03fc: douta_buf <= 22'h1000110101000100100110;
                12'h03fd: douta_buf <= 22'h0001010101100100100110;
                12'h03fe: douta_buf <= 22'h0101110110000100100110;
                12'h03ff: douta_buf <= 22'h1001110110000100100110;
                12'h0400: douta_buf <= 22'h0010010110100100100110;
                12'h0401: douta_buf <= 22'h0110110111000100100110;
                12'h0402: douta_buf <= 22'h1010110111000100100110;
                12'h0403: douta_buf <= 22'h0000001000011000000010;
                12'h0404: douta_buf <= 22'h0100101000111000000010;
                12'h0405: douta_buf <= 22'h1000101000111000000010;
                12'h0406: douta_buf <= 22'h0001001001011000000010;
                12'h0407: douta_buf <= 22'h0101101001111000000010;
                12'h0408: douta_buf <= 22'h1001101001111000000010;
                12'h0409: douta_buf <= 22'h0010001010011000000010;
                12'h040a: douta_buf <= 22'h0110101010111000000010;
                12'h040b: douta_buf <= 22'h1010101010111000000010;
                12'h040c: douta_buf <= 22'h0011001000001000000110;
                12'h040d: douta_buf <= 22'h0100011000101000100110;
                12'h040e: douta_buf <= 22'h1000011000101000100110;
                12'h040f: douta_buf <= 22'h0000111001001000100110;
                12'h0410: douta_buf <= 22'h0101011001101000100110;
                12'h0411: douta_buf <= 22'h1001011001101000100110;
                12'h0412: douta_buf <= 22'h0001111010001000100110;
                12'h0413: douta_buf <= 22'h0110011010101000100110;
                12'h0414: douta_buf <= 22'h1010011010101000100110;
                12'h0415: douta_buf <= 22'h0010111011001000100110;
                12'h0416: douta_buf <= 22'h0100001100011100000010;
                12'h0417: douta_buf <= 22'h1000001100011100000010;
                12'h0418: douta_buf <= 22'h0000101100111100000010;
                12'h0419: douta_buf <= 22'h0101001101011100000010;
                12'h041a: douta_buf <= 22'h1001001101011100000010;
                12'h041b: douta_buf <= 22'h0001101101111100000010;
                12'h041c: douta_buf <= 22'h0110001110011100000010;
                12'h041d: douta_buf <= 22'h1010001110011100000010;
                12'h041e: douta_buf <= 22'h0010101110111100000010;
                12'h041f: douta_buf <= 22'h0111001100001100000110;
                12'h0420: douta_buf <= 22'h1011001100001100000110;
                12'h0421: douta_buf <= 22'h0000011100101100100110;
                12'h0422: douta_buf <= 22'h0100111101001100100110;
                12'h0423: douta_buf <= 22'h1000111101001100100110;
                12'h0424: douta_buf <= 22'h0001011101101100100110;
                12'h0425: douta_buf <= 22'h0101111110001100100110;
                12'h0426: douta_buf <= 22'h1001111110001100100110;
                12'h0427: douta_buf <= 22'h0010011110101100100110;
                12'h0428: douta_buf <= 22'h0110111111001100100110;
                12'h0429: douta_buf <= 22'h1010111111001100100110;
                12'h042a: douta_buf <= 22'h0001101000000000000001;
                12'h042b: douta_buf <= 22'h0000000000000000000000;
                12'h042c: douta_buf <= 22'h0000000000000000000000;
                12'h042d: douta_buf <= 22'h0000000000000000000000;
                12'h042e: douta_buf <= 22'h0000000000000000000000;
                12'h042f: douta_buf <= 22'h0000000000010000000110;
                12'h0430: douta_buf <= 22'h0000100000110000000110;
                12'h0431: douta_buf <= 22'h0001000001010000000110;
                12'h0432: douta_buf <= 22'h0001100001110000000110;
                12'h0433: douta_buf <= 22'h0010000010010000000110;
                12'h0434: douta_buf <= 22'h0010100010110000000110;
                12'h0435: douta_buf <= 22'h0011000000000000000110;
                12'h0436: douta_buf <= 22'h0000010000100000000110;
                12'h0437: douta_buf <= 22'h0000110001000000000110;
                12'h0438: douta_buf <= 22'h0001010001100000000110;
                12'h0439: douta_buf <= 22'h0001110010000000000110;
                12'h043a: douta_buf <= 22'h0010010010100000000110;
                12'h043b: douta_buf <= 22'h0010110011000000000110;
                12'h043c: douta_buf <= 22'h0000000000010001001110;
                12'h043d: douta_buf <= 22'h0000100000110001001110;
                12'h043e: douta_buf <= 22'h0001000001010001001110;
                12'h043f: douta_buf <= 22'h0001100001110001001110;
                12'h0440: douta_buf <= 22'h0010000010010001001110;
                12'h0441: douta_buf <= 22'h0010100010110001001110;
                12'h0442: douta_buf <= 22'h0011000000000001001110;
                12'h0443: douta_buf <= 22'h0000010000100001001110;
                12'h0444: douta_buf <= 22'h0000110001000001001110;
                12'h0445: douta_buf <= 22'h0001010001100001001110;
                12'h0446: douta_buf <= 22'h0001110010000001001110;
                12'h0447: douta_buf <= 22'h0010010010100001001110;
                12'h0448: douta_buf <= 22'h0010110011000001001110;
                12'h0449: douta_buf <= 22'h0000000100010100000110;
                12'h044a: douta_buf <= 22'h0000100100110100000110;
                12'h044b: douta_buf <= 22'h0001000101010100000110;
                12'h044c: douta_buf <= 22'h0001100101110100000110;
                12'h044d: douta_buf <= 22'h0010000110010100000110;
                12'h044e: douta_buf <= 22'h0010100110110100000110;
                12'h044f: douta_buf <= 22'h0011000100000100000110;
                12'h0450: douta_buf <= 22'h0000010100100100000110;
                12'h0451: douta_buf <= 22'h0000110101000100000110;
                12'h0452: douta_buf <= 22'h0001010101100100000110;
                12'h0453: douta_buf <= 22'h0001110110000100000110;
                12'h0454: douta_buf <= 22'h0010010110100100000110;
                12'h0455: douta_buf <= 22'h0010110111000100000110;
                12'h0456: douta_buf <= 22'h0000000100010101001110;
                12'h0457: douta_buf <= 22'h0000100100110101001110;
                12'h0458: douta_buf <= 22'h0001000101010101001110;
                12'h0459: douta_buf <= 22'h0001100101110101001110;
                12'h045a: douta_buf <= 22'h0010000110010101001110;
                12'h045b: douta_buf <= 22'h0010100110110101001110;
                12'h045c: douta_buf <= 22'h0011000100000101001110;
                12'h045d: douta_buf <= 22'h0000010100100101001110;
                12'h045e: douta_buf <= 22'h0000110101000101001110;
                12'h045f: douta_buf <= 22'h0001010101100101001110;
                12'h0460: douta_buf <= 22'h0001110110000101001110;
                12'h0461: douta_buf <= 22'h0010010110100101001110;
                12'h0462: douta_buf <= 22'h0010110111000101001110;
                12'h0463: douta_buf <= 22'h0000001000011000000110;
                12'h0464: douta_buf <= 22'h0000101000111000000110;
                12'h0465: douta_buf <= 22'h0001001001011000000110;
                12'h0466: douta_buf <= 22'h0001101001111000000110;
                12'h0467: douta_buf <= 22'h0010001010011000000110;
                12'h0468: douta_buf <= 22'h0010101010111000000110;
                12'h0469: douta_buf <= 22'h0011001000001000000110;
                12'h046a: douta_buf <= 22'h0000011000101000000110;
                12'h046b: douta_buf <= 22'h0000111001001000000110;
                12'h046c: douta_buf <= 22'h0001011001101000000110;
                12'h046d: douta_buf <= 22'h0001111010001000000110;
                12'h046e: douta_buf <= 22'h0010011010101000000110;
                12'h046f: douta_buf <= 22'h0010111011001000000110;
                12'h0470: douta_buf <= 22'h0000001000011001001110;
                12'h0471: douta_buf <= 22'h0000101000111001001110;
                12'h0472: douta_buf <= 22'h0001001001011001001110;
                12'h0473: douta_buf <= 22'h0001101001111001001110;
                12'h0474: douta_buf <= 22'h0010001010011001001110;
                12'h0475: douta_buf <= 22'h0010101010111001001110;
                12'h0476: douta_buf <= 22'h0011001000001001001110;
                12'h0477: douta_buf <= 22'h0000011000101001001110;
                12'h0478: douta_buf <= 22'h0000111001001001001110;
                12'h0479: douta_buf <= 22'h0001011001101001001110;
                12'h047a: douta_buf <= 22'h0001111010001001001110;
                12'h047b: douta_buf <= 22'h0010011010101001001110;
                12'h047c: douta_buf <= 22'h0010111011001001001110;
                12'h047d: douta_buf <= 22'h0000001100011100000110;
                12'h047e: douta_buf <= 22'h0000101100111100000110;
                12'h047f: douta_buf <= 22'h0001001101011100000110;
                12'h0480: douta_buf <= 22'h0001101101111100000110;
                12'h0481: douta_buf <= 22'h0010001110011100000110;
                12'h0482: douta_buf <= 22'h0010101110111100000110;
                12'h0483: douta_buf <= 22'h0011001100001100000110;
                12'h0484: douta_buf <= 22'h0000011100101100000110;
                12'h0485: douta_buf <= 22'h0000111101001100000110;
                12'h0486: douta_buf <= 22'h0001011101101100000110;
                12'h0487: douta_buf <= 22'h0001111110001100000110;
                12'h0488: douta_buf <= 22'h0010011110101100000110;
                12'h0489: douta_buf <= 22'h0010111111001100000110;
                12'h048a: douta_buf <= 22'h0000001100011101001110;
                12'h048b: douta_buf <= 22'h0000101100111101001110;
                12'h048c: douta_buf <= 22'h0001001101011101001110;
                12'h048d: douta_buf <= 22'h0001101101111101001110;
                12'h048e: douta_buf <= 22'h0010001110011101001110;
                12'h048f: douta_buf <= 22'h0010101110111101001110;
                12'h0490: douta_buf <= 22'h0011001100001101001110;
                12'h0491: douta_buf <= 22'h0000011100101101001110;
                12'h0492: douta_buf <= 22'h0000111101001101001110;
                12'h0493: douta_buf <= 22'h0001011101101101001110;
                12'h0494: douta_buf <= 22'h0001111110001101001110;
                12'h0495: douta_buf <= 22'h0010011110101101001110;
                12'h0496: douta_buf <= 22'h0010111111001101001110;
                12'h0497: douta_buf <= 22'h0001101000000000000001;
                12'h0498: douta_buf <= 22'h0000000000000000000000;
                12'h0499: douta_buf <= 22'h0000000000000000000000;
                12'h049a: douta_buf <= 22'h0000000000000000000000;
                12'h049b: douta_buf <= 22'h0000000000000000000000;
                12'h049c: douta_buf <= 22'h0000000000010000000110;
                12'h049d: douta_buf <= 22'h0100100000110000000110;
                12'h049e: douta_buf <= 22'h1000100000110000000110;
                12'h049f: douta_buf <= 22'h0001000001010000000110;
                12'h04a0: douta_buf <= 22'h0101100001110000000110;
                12'h04a1: douta_buf <= 22'h1001100001110000000110;
                12'h04a2: douta_buf <= 22'h0010000010010000000110;
                12'h04a3: douta_buf <= 22'h0110100010110000000110;
                12'h04a4: douta_buf <= 22'h1010100010110000000110;
                12'h04a5: douta_buf <= 22'h0011000000000000000110;
                12'h04a6: douta_buf <= 22'h0100010000100000000110;
                12'h04a7: douta_buf <= 22'h1000010000100000000110;
                12'h04a8: douta_buf <= 22'h0000110001000000000110;
                12'h04a9: douta_buf <= 22'h0101010001100000000110;
                12'h04aa: douta_buf <= 22'h1001010001100000000110;
                12'h04ab: douta_buf <= 22'h0001110010000000000110;
                12'h04ac: douta_buf <= 22'h0110010010100000000110;
                12'h04ad: douta_buf <= 22'h1010010010100000000110;
                12'h04ae: douta_buf <= 22'h0010110011000000000110;
                12'h04af: douta_buf <= 22'h0100000000010001001110;
                12'h04b0: douta_buf <= 22'h1000000000010001001110;
                12'h04b1: douta_buf <= 22'h0000100000110001001110;
                12'h04b2: douta_buf <= 22'h0101000001010001001110;
                12'h04b3: douta_buf <= 22'h1001000001010001001110;
                12'h04b4: douta_buf <= 22'h0001100001110001001110;
                12'h04b5: douta_buf <= 22'h0110000010010001001110;
                12'h04b6: douta_buf <= 22'h1010000010010001001110;
                12'h04b7: douta_buf <= 22'h0010100010110001001110;
                12'h04b8: douta_buf <= 22'h0111000000000001001110;
                12'h04b9: douta_buf <= 22'h1011000000000001001110;
                12'h04ba: douta_buf <= 22'h0000010000100001001110;
                12'h04bb: douta_buf <= 22'h0100110001000001001110;
                12'h04bc: douta_buf <= 22'h1000110001000001001110;
                12'h04bd: douta_buf <= 22'h0001010001100001001110;
                12'h04be: douta_buf <= 22'h0101110010000001001110;
                12'h04bf: douta_buf <= 22'h1001110010000001001110;
                12'h04c0: douta_buf <= 22'h0010010010100001001110;
                12'h04c1: douta_buf <= 22'h0110110011000001001110;
                12'h04c2: douta_buf <= 22'h1010110011000001001110;
                12'h04c3: douta_buf <= 22'h0000000100010100000110;
                12'h04c4: douta_buf <= 22'h0100100100110100000110;
                12'h04c5: douta_buf <= 22'h1000100100110100000110;
                12'h04c6: douta_buf <= 22'h0001000101010100000110;
                12'h04c7: douta_buf <= 22'h0101100101110100000110;
                12'h04c8: douta_buf <= 22'h1001100101110100000110;
                12'h04c9: douta_buf <= 22'h0010000110010100000110;
                12'h04ca: douta_buf <= 22'h0110100110110100000110;
                12'h04cb: douta_buf <= 22'h1010100110110100000110;
                12'h04cc: douta_buf <= 22'h0011000100000100000110;
                12'h04cd: douta_buf <= 22'h0100010100100100000110;
                12'h04ce: douta_buf <= 22'h1000010100100100000110;
                12'h04cf: douta_buf <= 22'h0000110101000100000110;
                12'h04d0: douta_buf <= 22'h0101010101100100000110;
                12'h04d1: douta_buf <= 22'h1001010101100100000110;
                12'h04d2: douta_buf <= 22'h0001110110000100000110;
                12'h04d3: douta_buf <= 22'h0110010110100100000110;
                12'h04d4: douta_buf <= 22'h1010010110100100000110;
                12'h04d5: douta_buf <= 22'h0010110111000100000110;
                12'h04d6: douta_buf <= 22'h0100000100010101001110;
                12'h04d7: douta_buf <= 22'h1000000100010101001110;
                12'h04d8: douta_buf <= 22'h0000100100110101001110;
                12'h04d9: douta_buf <= 22'h0101000101010101001110;
                12'h04da: douta_buf <= 22'h1001000101010101001110;
                12'h04db: douta_buf <= 22'h0001100101110101001110;
                12'h04dc: douta_buf <= 22'h0110000110010101001110;
                12'h04dd: douta_buf <= 22'h1010000110010101001110;
                12'h04de: douta_buf <= 22'h0010100110110101001110;
                12'h04df: douta_buf <= 22'h0111000100000101001110;
                12'h04e0: douta_buf <= 22'h1011000100000101001110;
                12'h04e1: douta_buf <= 22'h0000010100100101001110;
                12'h04e2: douta_buf <= 22'h0100110101000101001110;
                12'h04e3: douta_buf <= 22'h1000110101000101001110;
                12'h04e4: douta_buf <= 22'h0001010101100101001110;
                12'h04e5: douta_buf <= 22'h0101110110000101001110;
                12'h04e6: douta_buf <= 22'h1001110110000101001110;
                12'h04e7: douta_buf <= 22'h0010010110100101001110;
                12'h04e8: douta_buf <= 22'h0110110111000101001110;
                12'h04e9: douta_buf <= 22'h1010110111000101001110;
                12'h04ea: douta_buf <= 22'h0000001000011000000110;
                12'h04eb: douta_buf <= 22'h0100101000111000000110;
                12'h04ec: douta_buf <= 22'h1000101000111000000110;
                12'h04ed: douta_buf <= 22'h0001001001011000000110;
                12'h04ee: douta_buf <= 22'h0101101001111000000110;
                12'h04ef: douta_buf <= 22'h1001101001111000000110;
                12'h04f0: douta_buf <= 22'h0010001010011000000110;
                12'h04f1: douta_buf <= 22'h0110101010111000000110;
                12'h04f2: douta_buf <= 22'h1010101010111000000110;
                12'h04f3: douta_buf <= 22'h0011001000001000000110;
                12'h04f4: douta_buf <= 22'h0100011000101000000110;
                12'h04f5: douta_buf <= 22'h1000011000101000000110;
                12'h04f6: douta_buf <= 22'h0000111001001000000110;
                12'h04f7: douta_buf <= 22'h0101011001101000000110;
                12'h04f8: douta_buf <= 22'h1001011001101000000110;
                12'h04f9: douta_buf <= 22'h0001111010001000000110;
                12'h04fa: douta_buf <= 22'h0110011010101000000110;
                12'h04fb: douta_buf <= 22'h1010011010101000000110;
                12'h04fc: douta_buf <= 22'h0010111011001000000110;
                12'h04fd: douta_buf <= 22'h0100001000011001001110;
                12'h04fe: douta_buf <= 22'h1000001000011001001110;
                12'h04ff: douta_buf <= 22'h0000101000111001001110;
                12'h0500: douta_buf <= 22'h0101001001011001001110;
                12'h0501: douta_buf <= 22'h1001001001011001001110;
                12'h0502: douta_buf <= 22'h0001101001111001001110;
                12'h0503: douta_buf <= 22'h0110001010011001001110;
                12'h0504: douta_buf <= 22'h1010001010011001001110;
                12'h0505: douta_buf <= 22'h0010101010111001001110;
                12'h0506: douta_buf <= 22'h0111001000001001001110;
                12'h0507: douta_buf <= 22'h1011001000001001001110;
                12'h0508: douta_buf <= 22'h0000011000101001001110;
                12'h0509: douta_buf <= 22'h0100111001001001001110;
                12'h050a: douta_buf <= 22'h1000111001001001001110;
                12'h050b: douta_buf <= 22'h0001011001101001001110;
                12'h050c: douta_buf <= 22'h0101111010001001001110;
                12'h050d: douta_buf <= 22'h1001111010001001001110;
                12'h050e: douta_buf <= 22'h0010011010101001001110;
                12'h050f: douta_buf <= 22'h0110111011001001001110;
                12'h0510: douta_buf <= 22'h1010111011001001001110;
                12'h0511: douta_buf <= 22'h0000001100011100000110;
                12'h0512: douta_buf <= 22'h0100101100111100000110;
                12'h0513: douta_buf <= 22'h1000101100111100000110;
                12'h0514: douta_buf <= 22'h0001001101011100000110;
                12'h0515: douta_buf <= 22'h0101101101111100000110;
                12'h0516: douta_buf <= 22'h1001101101111100000110;
                12'h0517: douta_buf <= 22'h0010001110011100000110;
                12'h0518: douta_buf <= 22'h0110101110111100000110;
                12'h0519: douta_buf <= 22'h1010101110111100000110;
                12'h051a: douta_buf <= 22'h0011001100001100000110;
                12'h051b: douta_buf <= 22'h0100011100101100000110;
                12'h051c: douta_buf <= 22'h1000011100101100000110;
                12'h051d: douta_buf <= 22'h0000111101001100000110;
                12'h051e: douta_buf <= 22'h0101011101101100000110;
                12'h051f: douta_buf <= 22'h1001011101101100000110;
                12'h0520: douta_buf <= 22'h0001111110001100000110;
                12'h0521: douta_buf <= 22'h0110011110101100000110;
                12'h0522: douta_buf <= 22'h1010011110101100000110;
                12'h0523: douta_buf <= 22'h0010111111001100000110;
                12'h0524: douta_buf <= 22'h0100001100011101001110;
                12'h0525: douta_buf <= 22'h1000001100011101001110;
                12'h0526: douta_buf <= 22'h0000101100111101001110;
                12'h0527: douta_buf <= 22'h0101001101011101001110;
                12'h0528: douta_buf <= 22'h1001001101011101001110;
                12'h0529: douta_buf <= 22'h0001101101111101001110;
                12'h052a: douta_buf <= 22'h0110001110011101001110;
                12'h052b: douta_buf <= 22'h1010001110011101001110;
                12'h052c: douta_buf <= 22'h0010101110111101001110;
                12'h052d: douta_buf <= 22'h0111001100001101001110;
                12'h052e: douta_buf <= 22'h1011001100001101001110;
                12'h052f: douta_buf <= 22'h0000011100101101001110;
                12'h0530: douta_buf <= 22'h0100111101001101001110;
                12'h0531: douta_buf <= 22'h1000111101001101001110;
                12'h0532: douta_buf <= 22'h0001011101101101001110;
                12'h0533: douta_buf <= 22'h0101111110001101001110;
                12'h0534: douta_buf <= 22'h1001111110001101001110;
                12'h0535: douta_buf <= 22'h0010011110101101001110;
                12'h0536: douta_buf <= 22'h0110111111001101001110;
                12'h0537: douta_buf <= 22'h1010111111001101001110;
                12'h0538: douta_buf <= 22'h0001101000000000000001;
                12'h0539: douta_buf <= 22'h0000000000000000000000;
                12'h053a: douta_buf <= 22'h0000000000000000000000;
                12'h053b: douta_buf <= 22'h0000000000000000000000;
                12'h053c: douta_buf <= 22'h0000000000000000000000;
                12'h053d: douta_buf <= 22'h0000000000010000001010;
                12'h053e: douta_buf <= 22'h0100100000110000100010;
                12'h053f: douta_buf <= 22'h0000110001000000001010;
                12'h0540: douta_buf <= 22'h0101010001100000100010;
                12'h0541: douta_buf <= 22'h0001100001110000001010;
                12'h0542: douta_buf <= 22'h0110000010010000100010;
                12'h0543: douta_buf <= 22'h0010010010100000001010;
                12'h0544: douta_buf <= 22'h0110110011000000100010;
                12'h0545: douta_buf <= 22'h0011000000000000000110;
                12'h0546: douta_buf <= 22'h0100010000100000001010;
                12'h0547: douta_buf <= 22'h0000100000110001000110;
                12'h0548: douta_buf <= 22'h0101000001010000001010;
                12'h0549: douta_buf <= 22'h0001010001100001000110;
                12'h054a: douta_buf <= 22'h0101110010000000001010;
                12'h054b: douta_buf <= 22'h0010000010010001000110;
                12'h054c: douta_buf <= 22'h0110100010110000001010;
                12'h054d: douta_buf <= 22'h0010110011000001000110;
                12'h054e: douta_buf <= 22'h0100000000010001000110;
                12'h054f: douta_buf <= 22'h0000010000100000100010;
                12'h0550: douta_buf <= 22'h0100110001000001000110;
                12'h0551: douta_buf <= 22'h0001000001010000100010;
                12'h0552: douta_buf <= 22'h0101100001110001000110;
                12'h0553: douta_buf <= 22'h0001110010000000100010;
                12'h0554: douta_buf <= 22'h0110010010100001000110;
                12'h0555: douta_buf <= 22'h0010100010110000100010;
                12'h0556: douta_buf <= 22'h0111000000000001001110;
                12'h0557: douta_buf <= 22'h0000000000010001110110;
                12'h0558: douta_buf <= 22'h0100100000110010001110;
                12'h0559: douta_buf <= 22'h0000110001000001110110;
                12'h055a: douta_buf <= 22'h0101010001100010001110;
                12'h055b: douta_buf <= 22'h0001100001110001110110;
                12'h055c: douta_buf <= 22'h0110000010010010001110;
                12'h055d: douta_buf <= 22'h0010010010100001110110;
                12'h055e: douta_buf <= 22'h0110110011000010001110;
                12'h055f: douta_buf <= 22'h0011000000000001110010;
                12'h0560: douta_buf <= 22'h0100010000100001110110;
                12'h0561: douta_buf <= 22'h0000100000110010110010;
                12'h0562: douta_buf <= 22'h0101000001010001110110;
                12'h0563: douta_buf <= 22'h0001010001100010110010;
                12'h0564: douta_buf <= 22'h0101110010000001110110;
                12'h0565: douta_buf <= 22'h0010000010010010110010;
                12'h0566: douta_buf <= 22'h0110100010110001110110;
                12'h0567: douta_buf <= 22'h0010110011000010110010;
                12'h0568: douta_buf <= 22'h0100000000010010110010;
                12'h0569: douta_buf <= 22'h0000010000100010001110;
                12'h056a: douta_buf <= 22'h0100110001000010110010;
                12'h056b: douta_buf <= 22'h0001000001010010001110;
                12'h056c: douta_buf <= 22'h0101100001110010110010;
                12'h056d: douta_buf <= 22'h0001110010000010001110;
                12'h056e: douta_buf <= 22'h0110010010100010110010;
                12'h056f: douta_buf <= 22'h0010100010110010001110;
                12'h0570: douta_buf <= 22'h0111000000000110100010;
                12'h0571: douta_buf <= 22'h0000000100010100001010;
                12'h0572: douta_buf <= 22'h0100100100110100100010;
                12'h0573: douta_buf <= 22'h0000110101000100001010;
                12'h0574: douta_buf <= 22'h0101010101100100100010;
                12'h0575: douta_buf <= 22'h0001100101110100001010;
                12'h0576: douta_buf <= 22'h0110000110010100100010;
                12'h0577: douta_buf <= 22'h0010010110100100001010;
                12'h0578: douta_buf <= 22'h0110110111000100100010;
                12'h0579: douta_buf <= 22'h0011000100000100000110;
                12'h057a: douta_buf <= 22'h0100010100100100001010;
                12'h057b: douta_buf <= 22'h0000100100110101000110;
                12'h057c: douta_buf <= 22'h0101000101010100001010;
                12'h057d: douta_buf <= 22'h0001010101100101000110;
                12'h057e: douta_buf <= 22'h0101110110000100001010;
                12'h057f: douta_buf <= 22'h0010000110010101000110;
                12'h0580: douta_buf <= 22'h0110100110110100001010;
                12'h0581: douta_buf <= 22'h0010110111000101000110;
                12'h0582: douta_buf <= 22'h0100000100010101000110;
                12'h0583: douta_buf <= 22'h0000010100100100100010;
                12'h0584: douta_buf <= 22'h0100110101000101000110;
                12'h0585: douta_buf <= 22'h0001000101010100100010;
                12'h0586: douta_buf <= 22'h0101100101110101000110;
                12'h0587: douta_buf <= 22'h0001110110000100100010;
                12'h0588: douta_buf <= 22'h0110010110100101000110;
                12'h0589: douta_buf <= 22'h0010100110110100100010;
                12'h058a: douta_buf <= 22'h0111000100000101001110;
                12'h058b: douta_buf <= 22'h0000000100010101110110;
                12'h058c: douta_buf <= 22'h0100100100110110001110;
                12'h058d: douta_buf <= 22'h0000110101000101110110;
                12'h058e: douta_buf <= 22'h0101010101100110001110;
                12'h058f: douta_buf <= 22'h0001100101110101110110;
                12'h0590: douta_buf <= 22'h0110000110010110001110;
                12'h0591: douta_buf <= 22'h0010010110100101110110;
                12'h0592: douta_buf <= 22'h0110110111000110001110;
                12'h0593: douta_buf <= 22'h0011000100000101110010;
                12'h0594: douta_buf <= 22'h0100010100100101110110;
                12'h0595: douta_buf <= 22'h0000100100110110110010;
                12'h0596: douta_buf <= 22'h0101000101010101110110;
                12'h0597: douta_buf <= 22'h0001010101100110110010;
                12'h0598: douta_buf <= 22'h0101110110000101110110;
                12'h0599: douta_buf <= 22'h0010000110010110110010;
                12'h059a: douta_buf <= 22'h0110100110110101110110;
                12'h059b: douta_buf <= 22'h0010110111000110110010;
                12'h059c: douta_buf <= 22'h0100000100010110110010;
                12'h059d: douta_buf <= 22'h0000010100100110001110;
                12'h059e: douta_buf <= 22'h0100110101000110110010;
                12'h059f: douta_buf <= 22'h0001000101010110001110;
                12'h05a0: douta_buf <= 22'h0101100101110110110010;
                12'h05a1: douta_buf <= 22'h0001110110000110001110;
                12'h05a2: douta_buf <= 22'h0110010110100110110010;
                12'h05a3: douta_buf <= 22'h0010100110110110001110;
                12'h05a4: douta_buf <= 22'h0111000100001010100010;
                12'h05a5: douta_buf <= 22'h0000001000011000001010;
                12'h05a6: douta_buf <= 22'h0100101000111000100010;
                12'h05a7: douta_buf <= 22'h0000111001001000001010;
                12'h05a8: douta_buf <= 22'h0101011001101000100010;
                12'h05a9: douta_buf <= 22'h0001101001111000001010;
                12'h05aa: douta_buf <= 22'h0110001010011000100010;
                12'h05ab: douta_buf <= 22'h0010011010101000001010;
                12'h05ac: douta_buf <= 22'h0110111011001000100010;
                12'h05ad: douta_buf <= 22'h0011001000001000000110;
                12'h05ae: douta_buf <= 22'h0100011000101000001010;
                12'h05af: douta_buf <= 22'h0000101000111001000110;
                12'h05b0: douta_buf <= 22'h0101001001011000001010;
                12'h05b1: douta_buf <= 22'h0001011001101001000110;
                12'h05b2: douta_buf <= 22'h0101111010001000001010;
                12'h05b3: douta_buf <= 22'h0010001010011001000110;
                12'h05b4: douta_buf <= 22'h0110101010111000001010;
                12'h05b5: douta_buf <= 22'h0010111011001001000110;
                12'h05b6: douta_buf <= 22'h0100001000011001000110;
                12'h05b7: douta_buf <= 22'h0000011000101000100010;
                12'h05b8: douta_buf <= 22'h0100111001001001000110;
                12'h05b9: douta_buf <= 22'h0001001001011000100010;
                12'h05ba: douta_buf <= 22'h0101101001111001000110;
                12'h05bb: douta_buf <= 22'h0001111010001000100010;
                12'h05bc: douta_buf <= 22'h0110011010101001000110;
                12'h05bd: douta_buf <= 22'h0010101010111000100010;
                12'h05be: douta_buf <= 22'h0111001000001001001110;
                12'h05bf: douta_buf <= 22'h0000001000011001110110;
                12'h05c0: douta_buf <= 22'h0100101000111010001110;
                12'h05c1: douta_buf <= 22'h0000111001001001110110;
                12'h05c2: douta_buf <= 22'h0101011001101010001110;
                12'h05c3: douta_buf <= 22'h0001101001111001110110;
                12'h05c4: douta_buf <= 22'h0110001010011010001110;
                12'h05c5: douta_buf <= 22'h0010011010101001110110;
                12'h05c6: douta_buf <= 22'h0110111011001010001110;
                12'h05c7: douta_buf <= 22'h0011001000001001110010;
                12'h05c8: douta_buf <= 22'h0100011000101001110110;
                12'h05c9: douta_buf <= 22'h0000101000111010110010;
                12'h05ca: douta_buf <= 22'h0101001001011001110110;
                12'h05cb: douta_buf <= 22'h0001011001101010110010;
                12'h05cc: douta_buf <= 22'h0101111010001001110110;
                12'h05cd: douta_buf <= 22'h0010001010011010110010;
                12'h05ce: douta_buf <= 22'h0110101010111001110110;
                12'h05cf: douta_buf <= 22'h0010111011001010110010;
                12'h05d0: douta_buf <= 22'h0100001000011010110010;
                12'h05d1: douta_buf <= 22'h0000011000101010001110;
                12'h05d2: douta_buf <= 22'h0100111001001010110010;
                12'h05d3: douta_buf <= 22'h0001001001011010001110;
                12'h05d4: douta_buf <= 22'h0101101001111010110010;
                12'h05d5: douta_buf <= 22'h0001111010001010001110;
                12'h05d6: douta_buf <= 22'h0110011010101010110010;
                12'h05d7: douta_buf <= 22'h0010101010111010001110;
                12'h05d8: douta_buf <= 22'h0111001000001110100010;
                12'h05d9: douta_buf <= 22'h0000001100011100001010;
                12'h05da: douta_buf <= 22'h0100101100111100100010;
                12'h05db: douta_buf <= 22'h0000111101001100001010;
                12'h05dc: douta_buf <= 22'h0101011101101100100010;
                12'h05dd: douta_buf <= 22'h0001101101111100001010;
                12'h05de: douta_buf <= 22'h0110001110011100100010;
                12'h05df: douta_buf <= 22'h0010011110101100001010;
                12'h05e0: douta_buf <= 22'h0110111111001100100010;
                12'h05e1: douta_buf <= 22'h0011001100001100000110;
                12'h05e2: douta_buf <= 22'h0100011100101100001010;
                12'h05e3: douta_buf <= 22'h0000101100111101000110;
                12'h05e4: douta_buf <= 22'h0101001101011100001010;
                12'h05e5: douta_buf <= 22'h0001011101101101000110;
                12'h05e6: douta_buf <= 22'h0101111110001100001010;
                12'h05e7: douta_buf <= 22'h0010001110011101000110;
                12'h05e8: douta_buf <= 22'h0110101110111100001010;
                12'h05e9: douta_buf <= 22'h0010111111001101000110;
                12'h05ea: douta_buf <= 22'h0100001100011101000110;
                12'h05eb: douta_buf <= 22'h0000011100101100100010;
                12'h05ec: douta_buf <= 22'h0100111101001101000110;
                12'h05ed: douta_buf <= 22'h0001001101011100100010;
                12'h05ee: douta_buf <= 22'h0101101101111101000110;
                12'h05ef: douta_buf <= 22'h0001111110001100100010;
                12'h05f0: douta_buf <= 22'h0110011110101101000110;
                12'h05f1: douta_buf <= 22'h0010101110111100100010;
                12'h05f2: douta_buf <= 22'h0111001100001101001110;
                12'h05f3: douta_buf <= 22'h0000001100011101110110;
                12'h05f4: douta_buf <= 22'h0100101100111110001110;
                12'h05f5: douta_buf <= 22'h0000111101001101110110;
                12'h05f6: douta_buf <= 22'h0101011101101110001110;
                12'h05f7: douta_buf <= 22'h0001101101111101110110;
                12'h05f8: douta_buf <= 22'h0110001110011110001110;
                12'h05f9: douta_buf <= 22'h0010011110101101110110;
                12'h05fa: douta_buf <= 22'h0110111111001110001110;
                12'h05fb: douta_buf <= 22'h0011001100001101110010;
                12'h05fc: douta_buf <= 22'h0100011100101101110110;
                12'h05fd: douta_buf <= 22'h0000101100111110110010;
                12'h05fe: douta_buf <= 22'h0101001101011101110110;
                12'h05ff: douta_buf <= 22'h0001011101101110110010;
                12'h0600: douta_buf <= 22'h0101111110001101110110;
                12'h0601: douta_buf <= 22'h0010001110011110110010;
                12'h0602: douta_buf <= 22'h0110101110111101110110;
                12'h0603: douta_buf <= 22'h0010111111001110110010;
                12'h0604: douta_buf <= 22'h0100001100011110110010;
                12'h0605: douta_buf <= 22'h0000011100101110001110;
                12'h0606: douta_buf <= 22'h0100111101001110110010;
                12'h0607: douta_buf <= 22'h0001001101011110001110;
                12'h0608: douta_buf <= 22'h0101101101111110110010;
                12'h0609: douta_buf <= 22'h0001111110001110001110;
                12'h060a: douta_buf <= 22'h0110011110101110110010;
                12'h060b: douta_buf <= 22'h0010101110111110001110;
                12'h060c: douta_buf <= 22'h0111001100000010100010;
                12'h060d: douta_buf <= 22'h0001101000000000000001;
                12'h060e: douta_buf <= 22'h0000000000000000000000;
                12'h060f: douta_buf <= 22'h0000000000000000000000;
                12'h0610: douta_buf <= 22'h0000000000000000000000;
                12'h0611: douta_buf <= 22'h0000000000000000000000;
                12'h0612: douta_buf <= 22'h0000000000010000001010;
                12'h0613: douta_buf <= 22'h0100100000110000100010;
                12'h0614: douta_buf <= 22'h1000100000110000100010;
                12'h0615: douta_buf <= 22'h0001000001010001000110;
                12'h0616: douta_buf <= 22'h0101100001110000001010;
                12'h0617: douta_buf <= 22'h1001100001110000001010;
                12'h0618: douta_buf <= 22'h0010000010010000100010;
                12'h0619: douta_buf <= 22'h0110100010110001000110;
                12'h061a: douta_buf <= 22'h1010100010110001000110;
                12'h061b: douta_buf <= 22'h0011000000000000000110;
                12'h061c: douta_buf <= 22'h0100010000100000001010;
                12'h061d: douta_buf <= 22'h1000010000100000001010;
                12'h061e: douta_buf <= 22'h0000110001000000100010;
                12'h061f: douta_buf <= 22'h0101010001100001000110;
                12'h0620: douta_buf <= 22'h1001010001100001000110;
                12'h0621: douta_buf <= 22'h0001110010000000001010;
                12'h0622: douta_buf <= 22'h0110010010100000100010;
                12'h0623: douta_buf <= 22'h1010010010100000100010;
                12'h0624: douta_buf <= 22'h0010110011000001000110;
                12'h0625: douta_buf <= 22'h0100000000010001000110;
                12'h0626: douta_buf <= 22'h1000000000010001000110;
                12'h0627: douta_buf <= 22'h0000100000110000001010;
                12'h0628: douta_buf <= 22'h0101000001010000100010;
                12'h0629: douta_buf <= 22'h1001000001010000100010;
                12'h062a: douta_buf <= 22'h0001100001110001000110;
                12'h062b: douta_buf <= 22'h0110000010010000001010;
                12'h062c: douta_buf <= 22'h1010000010010000001010;
                12'h062d: douta_buf <= 22'h0010100010110000100010;
                12'h062e: douta_buf <= 22'h0111000000000001001110;
                12'h062f: douta_buf <= 22'h1011000000000001001110;
                12'h0630: douta_buf <= 22'h0000010000100010110010;
                12'h0631: douta_buf <= 22'h0100110001000001110110;
                12'h0632: douta_buf <= 22'h1000110001000001110110;
                12'h0633: douta_buf <= 22'h0001010001100010001110;
                12'h0634: douta_buf <= 22'h0101110010000010110010;
                12'h0635: douta_buf <= 22'h1001110010000010110010;
                12'h0636: douta_buf <= 22'h0010010010100001110110;
                12'h0637: douta_buf <= 22'h0110110011000010001110;
                12'h0638: douta_buf <= 22'h1010110011000010001110;
                12'h0639: douta_buf <= 22'h0000000000010010001110;
                12'h063a: douta_buf <= 22'h0100100000110010110010;
                12'h063b: douta_buf <= 22'h1000100000110010110010;
                12'h063c: douta_buf <= 22'h0001000001010001110110;
                12'h063d: douta_buf <= 22'h0101100001110010001110;
                12'h063e: douta_buf <= 22'h1001100001110010001110;
                12'h063f: douta_buf <= 22'h0010000010010010110010;
                12'h0640: douta_buf <= 22'h0110100010110001110110;
                12'h0641: douta_buf <= 22'h1010100010110001110110;
                12'h0642: douta_buf <= 22'h0011000000000010010110;
                12'h0643: douta_buf <= 22'h0100010000100010001110;
                12'h0644: douta_buf <= 22'h1000010000100010001110;
                12'h0645: douta_buf <= 22'h0000110001000010110010;
                12'h0646: douta_buf <= 22'h0101010001100001110110;
                12'h0647: douta_buf <= 22'h1001010001100001110110;
                12'h0648: douta_buf <= 22'h0001110010000010001110;
                12'h0649: douta_buf <= 22'h0110010010100010110010;
                12'h064a: douta_buf <= 22'h1010010010100010110010;
                12'h064b: douta_buf <= 22'h0010110011000001110110;
                12'h064c: douta_buf <= 22'h0100000100010100001010;
                12'h064d: douta_buf <= 22'h1000000100010100001010;
                12'h064e: douta_buf <= 22'h0000100100110100100010;
                12'h064f: douta_buf <= 22'h0101000101010101000110;
                12'h0650: douta_buf <= 22'h1001000101010101000110;
                12'h0651: douta_buf <= 22'h0001100101110100001010;
                12'h0652: douta_buf <= 22'h0110000110010100100010;
                12'h0653: douta_buf <= 22'h1010000110010100100010;
                12'h0654: douta_buf <= 22'h0010100110110101000110;
                12'h0655: douta_buf <= 22'h0111000100000100000110;
                12'h0656: douta_buf <= 22'h1011000100000100000110;
                12'h0657: douta_buf <= 22'h0000010100100100001010;
                12'h0658: douta_buf <= 22'h0100110101000100100010;
                12'h0659: douta_buf <= 22'h1000110101000100100010;
                12'h065a: douta_buf <= 22'h0001010101100101000110;
                12'h065b: douta_buf <= 22'h0101110110000100001010;
                12'h065c: douta_buf <= 22'h1001110110000100001010;
                12'h065d: douta_buf <= 22'h0010010110100100100010;
                12'h065e: douta_buf <= 22'h0110110111000101000110;
                12'h065f: douta_buf <= 22'h1010110111000101000110;
                12'h0660: douta_buf <= 22'h0000000100010101000110;
                12'h0661: douta_buf <= 22'h0100100100110100001010;
                12'h0662: douta_buf <= 22'h1000100100110100001010;
                12'h0663: douta_buf <= 22'h0001000101010100100010;
                12'h0664: douta_buf <= 22'h0101100101110101000110;
                12'h0665: douta_buf <= 22'h1001100101110101000110;
                12'h0666: douta_buf <= 22'h0010000110010100001010;
                12'h0667: douta_buf <= 22'h0110100110110100100010;
                12'h0668: douta_buf <= 22'h1010100110110100100010;
                12'h0669: douta_buf <= 22'h0011000100000101001110;
                12'h066a: douta_buf <= 22'h0100010100100110110010;
                12'h066b: douta_buf <= 22'h1000010100100110110010;
                12'h066c: douta_buf <= 22'h0000110101000101110110;
                12'h066d: douta_buf <= 22'h0101010101100110001110;
                12'h066e: douta_buf <= 22'h1001010101100110001110;
                12'h066f: douta_buf <= 22'h0001110110000110110010;
                12'h0670: douta_buf <= 22'h0110010110100101110110;
                12'h0671: douta_buf <= 22'h1010010110100101110110;
                12'h0672: douta_buf <= 22'h0010110111000110001110;
                12'h0673: douta_buf <= 22'h0100000100010110001110;
                12'h0674: douta_buf <= 22'h1000000100010110001110;
                12'h0675: douta_buf <= 22'h0000100100110110110010;
                12'h0676: douta_buf <= 22'h0101000101010101110110;
                12'h0677: douta_buf <= 22'h1001000101010101110110;
                12'h0678: douta_buf <= 22'h0001100101110110001110;
                12'h0679: douta_buf <= 22'h0110000110010110110010;
                12'h067a: douta_buf <= 22'h1010000110010110110010;
                12'h067b: douta_buf <= 22'h0010100110110101110110;
                12'h067c: douta_buf <= 22'h0111000100000110010110;
                12'h067d: douta_buf <= 22'h1011000100000110010110;
                12'h067e: douta_buf <= 22'h0000010100100110001110;
                12'h067f: douta_buf <= 22'h0100110101000110110010;
                12'h0680: douta_buf <= 22'h1000110101000110110010;
                12'h0681: douta_buf <= 22'h0001010101100101110110;
                12'h0682: douta_buf <= 22'h0101110110000110001110;
                12'h0683: douta_buf <= 22'h1001110110000110001110;
                12'h0684: douta_buf <= 22'h0010010110100110110010;
                12'h0685: douta_buf <= 22'h0110110111000101110110;
                12'h0686: douta_buf <= 22'h1010110111000101110110;
                12'h0687: douta_buf <= 22'h0000001000011000001010;
                12'h0688: douta_buf <= 22'h0100101000111000100010;
                12'h0689: douta_buf <= 22'h1000101000111000100010;
                12'h068a: douta_buf <= 22'h0001001001011001000110;
                12'h068b: douta_buf <= 22'h0101101001111000001010;
                12'h068c: douta_buf <= 22'h1001101001111000001010;
                12'h068d: douta_buf <= 22'h0010001010011000100010;
                12'h068e: douta_buf <= 22'h0110101010111001000110;
                12'h068f: douta_buf <= 22'h1010101010111001000110;
                12'h0690: douta_buf <= 22'h0011001000001000000110;
                12'h0691: douta_buf <= 22'h0100011000101000001010;
                12'h0692: douta_buf <= 22'h1000011000101000001010;
                12'h0693: douta_buf <= 22'h0000111001001000100010;
                12'h0694: douta_buf <= 22'h0101011001101001000110;
                12'h0695: douta_buf <= 22'h1001011001101001000110;
                12'h0696: douta_buf <= 22'h0001111010001000001010;
                12'h0697: douta_buf <= 22'h0110011010101000100010;
                12'h0698: douta_buf <= 22'h1010011010101000100010;
                12'h0699: douta_buf <= 22'h0010111011001001000110;
                12'h069a: douta_buf <= 22'h0100001000011001000110;
                12'h069b: douta_buf <= 22'h1000001000011001000110;
                12'h069c: douta_buf <= 22'h0000101000111000001010;
                12'h069d: douta_buf <= 22'h0101001001011000100010;
                12'h069e: douta_buf <= 22'h1001001001011000100010;
                12'h069f: douta_buf <= 22'h0001101001111001000110;
                12'h06a0: douta_buf <= 22'h0110001010011000001010;
                12'h06a1: douta_buf <= 22'h1010001010011000001010;
                12'h06a2: douta_buf <= 22'h0010101010111000100010;
                12'h06a3: douta_buf <= 22'h0111001000001001001110;
                12'h06a4: douta_buf <= 22'h1011001000001001001110;
                12'h06a5: douta_buf <= 22'h0000011000101010110010;
                12'h06a6: douta_buf <= 22'h0100111001001001110110;
                12'h06a7: douta_buf <= 22'h1000111001001001110110;
                12'h06a8: douta_buf <= 22'h0001011001101010001110;
                12'h06a9: douta_buf <= 22'h0101111010001010110010;
                12'h06aa: douta_buf <= 22'h1001111010001010110010;
                12'h06ab: douta_buf <= 22'h0010011010101001110110;
                12'h06ac: douta_buf <= 22'h0110111011001010001110;
                12'h06ad: douta_buf <= 22'h1010111011001010001110;
                12'h06ae: douta_buf <= 22'h0000001000011010001110;
                12'h06af: douta_buf <= 22'h0100101000111010110010;
                12'h06b0: douta_buf <= 22'h1000101000111010110010;
                12'h06b1: douta_buf <= 22'h0001001001011001110110;
                12'h06b2: douta_buf <= 22'h0101101001111010001110;
                12'h06b3: douta_buf <= 22'h1001101001111010001110;
                12'h06b4: douta_buf <= 22'h0010001010011010110010;
                12'h06b5: douta_buf <= 22'h0110101010111001110110;
                12'h06b6: douta_buf <= 22'h1010101010111001110110;
                12'h06b7: douta_buf <= 22'h0011001000001010010110;
                12'h06b8: douta_buf <= 22'h0100011000101010001110;
                12'h06b9: douta_buf <= 22'h1000011000101010001110;
                12'h06ba: douta_buf <= 22'h0000111001001010110010;
                12'h06bb: douta_buf <= 22'h0101011001101001110110;
                12'h06bc: douta_buf <= 22'h1001011001101001110110;
                12'h06bd: douta_buf <= 22'h0001111010001010001110;
                12'h06be: douta_buf <= 22'h0110011010101010110010;
                12'h06bf: douta_buf <= 22'h1010011010101010110010;
                12'h06c0: douta_buf <= 22'h0010111011001001110110;
                12'h06c1: douta_buf <= 22'h0100001100011100001010;
                12'h06c2: douta_buf <= 22'h1000001100011100001010;
                12'h06c3: douta_buf <= 22'h0000101100111100100010;
                12'h06c4: douta_buf <= 22'h0101001101011101000110;
                12'h06c5: douta_buf <= 22'h1001001101011101000110;
                12'h06c6: douta_buf <= 22'h0001101101111100001010;
                12'h06c7: douta_buf <= 22'h0110001110011100100010;
                12'h06c8: douta_buf <= 22'h1010001110011100100010;
                12'h06c9: douta_buf <= 22'h0010101110111101000110;
                12'h06ca: douta_buf <= 22'h0111001100001100000110;
                12'h06cb: douta_buf <= 22'h1011001100001100000110;
                12'h06cc: douta_buf <= 22'h0000011100101100001010;
                12'h06cd: douta_buf <= 22'h0100111101001100100010;
                12'h06ce: douta_buf <= 22'h1000111101001100100010;
                12'h06cf: douta_buf <= 22'h0001011101101101000110;
                12'h06d0: douta_buf <= 22'h0101111110001100001010;
                12'h06d1: douta_buf <= 22'h1001111110001100001010;
                12'h06d2: douta_buf <= 22'h0010011110101100100010;
                12'h06d3: douta_buf <= 22'h0110111111001101000110;
                12'h06d4: douta_buf <= 22'h1010111111001101000110;
                12'h06d5: douta_buf <= 22'h0000001100011101000110;
                12'h06d6: douta_buf <= 22'h0100101100111100001010;
                12'h06d7: douta_buf <= 22'h1000101100111100001010;
                12'h06d8: douta_buf <= 22'h0001001101011100100010;
                12'h06d9: douta_buf <= 22'h0101101101111101000110;
                12'h06da: douta_buf <= 22'h1001101101111101000110;
                12'h06db: douta_buf <= 22'h0010001110011100001010;
                12'h06dc: douta_buf <= 22'h0110101110111100100010;
                12'h06dd: douta_buf <= 22'h1010101110111100100010;
                12'h06de: douta_buf <= 22'h0011001100001101001110;
                12'h06df: douta_buf <= 22'h0100011100101110110010;
                12'h06e0: douta_buf <= 22'h1000011100101110110010;
                12'h06e1: douta_buf <= 22'h0000111101001101110110;
                12'h06e2: douta_buf <= 22'h0101011101101110001110;
                12'h06e3: douta_buf <= 22'h1001011101101110001110;
                12'h06e4: douta_buf <= 22'h0001111110001110110010;
                12'h06e5: douta_buf <= 22'h0110011110101101110110;
                12'h06e6: douta_buf <= 22'h1010011110101101110110;
                12'h06e7: douta_buf <= 22'h0010111111001110001110;
                12'h06e8: douta_buf <= 22'h0100001100011110001110;
                12'h06e9: douta_buf <= 22'h1000001100011110001110;
                12'h06ea: douta_buf <= 22'h0000101100111110110010;
                12'h06eb: douta_buf <= 22'h0101001101011101110110;
                12'h06ec: douta_buf <= 22'h1001001101011101110110;
                12'h06ed: douta_buf <= 22'h0001101101111110001110;
                12'h06ee: douta_buf <= 22'h0110001110011110110010;
                12'h06ef: douta_buf <= 22'h1010001110011110110010;
                12'h06f0: douta_buf <= 22'h0010101110111101110110;
                12'h06f1: douta_buf <= 22'h0111001100001110010110;
                12'h06f2: douta_buf <= 22'h1011001100001110010110;
                12'h06f3: douta_buf <= 22'h0000011100101110001110;
                12'h06f4: douta_buf <= 22'h0100111101001110110010;
                12'h06f5: douta_buf <= 22'h1000111101001110110010;
                12'h06f6: douta_buf <= 22'h0001011101101101110110;
                12'h06f7: douta_buf <= 22'h0101111110001110001110;
                12'h06f8: douta_buf <= 22'h1001111110001110001110;
                12'h06f9: douta_buf <= 22'h0010011110101110110010;
                12'h06fa: douta_buf <= 22'h0110111111001101110110;
                12'h06fb: douta_buf <= 22'h1010111111001101110110;
                12'h06fc: douta_buf <= 22'h0001101000000000000001;
                12'h06fd: douta_buf <= 22'h0000000000000000000000;
                12'h06fe: douta_buf <= 22'h0000000000000000000000;
                12'h06ff: douta_buf <= 22'h0000000000000000000000;
                12'h0700: douta_buf <= 22'h0000000000000000000000;
                12'h0701: douta_buf <= 22'h0000000000010000001010;
                12'h0702: douta_buf <= 22'h0100100000110000100010;
                12'h0703: douta_buf <= 22'h1000100000110000100010;
                12'h0704: douta_buf <= 22'h0101000001010001000110;
                12'h0705: douta_buf <= 22'h1001000001010001000110;
                12'h0706: douta_buf <= 22'h0001100001110000001010;
                12'h0707: douta_buf <= 22'h0110000010010000100010;
                12'h0708: douta_buf <= 22'h1010000010010000100010;
                12'h0709: douta_buf <= 22'h0110100010110001000110;
                12'h070a: douta_buf <= 22'h1010100010110001000110;
                12'h070b: douta_buf <= 22'h0011000000000000000110;
                12'h070c: douta_buf <= 22'h0100010000100000001010;
                12'h070d: douta_buf <= 22'h1000010000100000001010;
                12'h070e: douta_buf <= 22'h0100110001000000100010;
                12'h070f: douta_buf <= 22'h1000110001000000100010;
                12'h0710: douta_buf <= 22'h0001010001100001000110;
                12'h0711: douta_buf <= 22'h0101110010000000001010;
                12'h0712: douta_buf <= 22'h1001110010000000001010;
                12'h0713: douta_buf <= 22'h0110010010100000100010;
                12'h0714: douta_buf <= 22'h1010010010100000100010;
                12'h0715: douta_buf <= 22'h0010110011000001000110;
                12'h0716: douta_buf <= 22'h0100000000010001000110;
                12'h0717: douta_buf <= 22'h1000000000010001000110;
                12'h0718: douta_buf <= 22'h0100100000110000001010;
                12'h0719: douta_buf <= 22'h1000100000110000001010;
                12'h071a: douta_buf <= 22'h0001000001010000100010;
                12'h071b: douta_buf <= 22'h0101100001110001000110;
                12'h071c: douta_buf <= 22'h1001100001110001000110;
                12'h071d: douta_buf <= 22'h0110000010010000001010;
                12'h071e: douta_buf <= 22'h1010000010010000001010;
                12'h071f: douta_buf <= 22'h0010100010110000100010;
                12'h0720: douta_buf <= 22'h0111000000000001001110;
                12'h0721: douta_buf <= 22'h1011000000000001001110;
                12'h0722: douta_buf <= 22'h0100010000100010110010;
                12'h0723: douta_buf <= 22'h1000010000100010110010;
                12'h0724: douta_buf <= 22'h0000110001000001110110;
                12'h0725: douta_buf <= 22'h0101010001100010001110;
                12'h0726: douta_buf <= 22'h1001010001100010001110;
                12'h0727: douta_buf <= 22'h0101110010000010110010;
                12'h0728: douta_buf <= 22'h1001110010000010110010;
                12'h0729: douta_buf <= 22'h0010010010100001110110;
                12'h072a: douta_buf <= 22'h0110110011000010001110;
                12'h072b: douta_buf <= 22'h1010110011000010001110;
                12'h072c: douta_buf <= 22'h0100000000010010001110;
                12'h072d: douta_buf <= 22'h1000000000010010001110;
                12'h072e: douta_buf <= 22'h0000100000110010110010;
                12'h072f: douta_buf <= 22'h0101000001010001110110;
                12'h0730: douta_buf <= 22'h1001000001010001110110;
                12'h0731: douta_buf <= 22'h0101100001110010001110;
                12'h0732: douta_buf <= 22'h1001100001110010001110;
                12'h0733: douta_buf <= 22'h0010000010010010110010;
                12'h0734: douta_buf <= 22'h0110100010110001110110;
                12'h0735: douta_buf <= 22'h1010100010110001110110;
                12'h0736: douta_buf <= 22'h0111000000000010010110;
                12'h0737: douta_buf <= 22'h1011000000000010010110;
                12'h0738: douta_buf <= 22'h0000010000100010001110;
                12'h0739: douta_buf <= 22'h0100110001000010110010;
                12'h073a: douta_buf <= 22'h1000110001000010110010;
                12'h073b: douta_buf <= 22'h0101010001100001110110;
                12'h073c: douta_buf <= 22'h1001010001100001110110;
                12'h073d: douta_buf <= 22'h0001110010000010001110;
                12'h073e: douta_buf <= 22'h0110010010100010110010;
                12'h073f: douta_buf <= 22'h1010010010100010110010;
                12'h0740: douta_buf <= 22'h0110110011000001110110;
                12'h0741: douta_buf <= 22'h1010110011000001110110;
                12'h0742: douta_buf <= 22'h0000000100010100001010;
                12'h0743: douta_buf <= 22'h0100100100110100100010;
                12'h0744: douta_buf <= 22'h1000100100110100100010;
                12'h0745: douta_buf <= 22'h0101000101010101000110;
                12'h0746: douta_buf <= 22'h1001000101010101000110;
                12'h0747: douta_buf <= 22'h0001100101110100001010;
                12'h0748: douta_buf <= 22'h0110000110010100100010;
                12'h0749: douta_buf <= 22'h1010000110010100100010;
                12'h074a: douta_buf <= 22'h0110100110110101000110;
                12'h074b: douta_buf <= 22'h1010100110110101000110;
                12'h074c: douta_buf <= 22'h0011000100000100000110;
                12'h074d: douta_buf <= 22'h0100010100100100001010;
                12'h074e: douta_buf <= 22'h1000010100100100001010;
                12'h074f: douta_buf <= 22'h0100110101000100100010;
                12'h0750: douta_buf <= 22'h1000110101000100100010;
                12'h0751: douta_buf <= 22'h0001010101100101000110;
                12'h0752: douta_buf <= 22'h0101110110000100001010;
                12'h0753: douta_buf <= 22'h1001110110000100001010;
                12'h0754: douta_buf <= 22'h0110010110100100100010;
                12'h0755: douta_buf <= 22'h1010010110100100100010;
                12'h0756: douta_buf <= 22'h0010110111000101000110;
                12'h0757: douta_buf <= 22'h0100000100010101000110;
                12'h0758: douta_buf <= 22'h1000000100010101000110;
                12'h0759: douta_buf <= 22'h0100100100110100001010;
                12'h075a: douta_buf <= 22'h1000100100110100001010;
                12'h075b: douta_buf <= 22'h0001000101010100100010;
                12'h075c: douta_buf <= 22'h0101100101110101000110;
                12'h075d: douta_buf <= 22'h1001100101110101000110;
                12'h075e: douta_buf <= 22'h0110000110010100001010;
                12'h075f: douta_buf <= 22'h1010000110010100001010;
                12'h0760: douta_buf <= 22'h0010100110110100100010;
                12'h0761: douta_buf <= 22'h0111000100000101001110;
                12'h0762: douta_buf <= 22'h1011000100000101001110;
                12'h0763: douta_buf <= 22'h0100010100100110110010;
                12'h0764: douta_buf <= 22'h1000010100100110110010;
                12'h0765: douta_buf <= 22'h0000110101000101110110;
                12'h0766: douta_buf <= 22'h0101010101100110001110;
                12'h0767: douta_buf <= 22'h1001010101100110001110;
                12'h0768: douta_buf <= 22'h0101110110000110110010;
                12'h0769: douta_buf <= 22'h1001110110000110110010;
                12'h076a: douta_buf <= 22'h0010010110100101110110;
                12'h076b: douta_buf <= 22'h0110110111000110001110;
                12'h076c: douta_buf <= 22'h1010110111000110001110;
                12'h076d: douta_buf <= 22'h0100000100010110001110;
                12'h076e: douta_buf <= 22'h1000000100010110001110;
                12'h076f: douta_buf <= 22'h0000100100110110110010;
                12'h0770: douta_buf <= 22'h0101000101010101110110;
                12'h0771: douta_buf <= 22'h1001000101010101110110;
                12'h0772: douta_buf <= 22'h0101100101110110001110;
                12'h0773: douta_buf <= 22'h1001100101110110001110;
                12'h0774: douta_buf <= 22'h0010000110010110110010;
                12'h0775: douta_buf <= 22'h0110100110110101110110;
                12'h0776: douta_buf <= 22'h1010100110110101110110;
                12'h0777: douta_buf <= 22'h0111000100000110010110;
                12'h0778: douta_buf <= 22'h1011000100000110010110;
                12'h0779: douta_buf <= 22'h0000010100100110001110;
                12'h077a: douta_buf <= 22'h0100110101000110110010;
                12'h077b: douta_buf <= 22'h1000110101000110110010;
                12'h077c: douta_buf <= 22'h0101010101100101110110;
                12'h077d: douta_buf <= 22'h1001010101100101110110;
                12'h077e: douta_buf <= 22'h0001110110000110001110;
                12'h077f: douta_buf <= 22'h0110010110100110110010;
                12'h0780: douta_buf <= 22'h1010010110100110110010;
                12'h0781: douta_buf <= 22'h0110110111000101110110;
                12'h0782: douta_buf <= 22'h1010110111000101110110;
                12'h0783: douta_buf <= 22'h0000001000011000001010;
                12'h0784: douta_buf <= 22'h0100101000111000100010;
                12'h0785: douta_buf <= 22'h1000101000111000100010;
                12'h0786: douta_buf <= 22'h0101001001011001000110;
                12'h0787: douta_buf <= 22'h1001001001011001000110;
                12'h0788: douta_buf <= 22'h0001101001111000001010;
                12'h0789: douta_buf <= 22'h0110001010011000100010;
                12'h078a: douta_buf <= 22'h1010001010011000100010;
                12'h078b: douta_buf <= 22'h0110101010111001000110;
                12'h078c: douta_buf <= 22'h1010101010111001000110;
                12'h078d: douta_buf <= 22'h0011001000001000000110;
                12'h078e: douta_buf <= 22'h0100011000101000001010;
                12'h078f: douta_buf <= 22'h1000011000101000001010;
                12'h0790: douta_buf <= 22'h0100111001001000100010;
                12'h0791: douta_buf <= 22'h1000111001001000100010;
                12'h0792: douta_buf <= 22'h0001011001101001000110;
                12'h0793: douta_buf <= 22'h0101111010001000001010;
                12'h0794: douta_buf <= 22'h1001111010001000001010;
                12'h0795: douta_buf <= 22'h0110011010101000100010;
                12'h0796: douta_buf <= 22'h1010011010101000100010;
                12'h0797: douta_buf <= 22'h0010111011001001000110;
                12'h0798: douta_buf <= 22'h0100001000011001000110;
                12'h0799: douta_buf <= 22'h1000001000011001000110;
                12'h079a: douta_buf <= 22'h0100101000111000001010;
                12'h079b: douta_buf <= 22'h1000101000111000001010;
                12'h079c: douta_buf <= 22'h0001001001011000100010;
                12'h079d: douta_buf <= 22'h0101101001111001000110;
                12'h079e: douta_buf <= 22'h1001101001111001000110;
                12'h079f: douta_buf <= 22'h0110001010011000001010;
                12'h07a0: douta_buf <= 22'h1010001010011000001010;
                12'h07a1: douta_buf <= 22'h0010101010111000100010;
                12'h07a2: douta_buf <= 22'h0111001000001001001110;
                12'h07a3: douta_buf <= 22'h1011001000001001001110;
                12'h07a4: douta_buf <= 22'h0100011000101010110010;
                12'h07a5: douta_buf <= 22'h1000011000101010110010;
                12'h07a6: douta_buf <= 22'h0000111001001001110110;
                12'h07a7: douta_buf <= 22'h0101011001101010001110;
                12'h07a8: douta_buf <= 22'h1001011001101010001110;
                12'h07a9: douta_buf <= 22'h0101111010001010110010;
                12'h07aa: douta_buf <= 22'h1001111010001010110010;
                12'h07ab: douta_buf <= 22'h0010011010101001110110;
                12'h07ac: douta_buf <= 22'h0110111011001010001110;
                12'h07ad: douta_buf <= 22'h1010111011001010001110;
                12'h07ae: douta_buf <= 22'h0100001000011010001110;
                12'h07af: douta_buf <= 22'h1000001000011010001110;
                12'h07b0: douta_buf <= 22'h0000101000111010110010;
                12'h07b1: douta_buf <= 22'h0101001001011001110110;
                12'h07b2: douta_buf <= 22'h1001001001011001110110;
                12'h07b3: douta_buf <= 22'h0101101001111010001110;
                12'h07b4: douta_buf <= 22'h1001101001111010001110;
                12'h07b5: douta_buf <= 22'h0010001010011010110010;
                12'h07b6: douta_buf <= 22'h0110101010111001110110;
                12'h07b7: douta_buf <= 22'h1010101010111001110110;
                12'h07b8: douta_buf <= 22'h0111001000001010010110;
                12'h07b9: douta_buf <= 22'h1011001000001010010110;
                12'h07ba: douta_buf <= 22'h0000011000101010001110;
                12'h07bb: douta_buf <= 22'h0100111001001010110010;
                12'h07bc: douta_buf <= 22'h1000111001001010110010;
                12'h07bd: douta_buf <= 22'h0101011001101001110110;
                12'h07be: douta_buf <= 22'h1001011001101001110110;
                12'h07bf: douta_buf <= 22'h0001111010001010001110;
                12'h07c0: douta_buf <= 22'h0110011010101010110010;
                12'h07c1: douta_buf <= 22'h1010011010101010110010;
                12'h07c2: douta_buf <= 22'h0110111011001001110110;
                12'h07c3: douta_buf <= 22'h1010111011001001110110;
                12'h07c4: douta_buf <= 22'h0000001100011100001010;
                12'h07c5: douta_buf <= 22'h0100101100111100100010;
                12'h07c6: douta_buf <= 22'h1000101100111100100010;
                12'h07c7: douta_buf <= 22'h0101001101011101000110;
                12'h07c8: douta_buf <= 22'h1001001101011101000110;
                12'h07c9: douta_buf <= 22'h0001101101111100001010;
                12'h07ca: douta_buf <= 22'h0110001110011100100010;
                12'h07cb: douta_buf <= 22'h1010001110011100100010;
                12'h07cc: douta_buf <= 22'h0110101110111101000110;
                12'h07cd: douta_buf <= 22'h1010101110111101000110;
                12'h07ce: douta_buf <= 22'h0011001100001100000110;
                12'h07cf: douta_buf <= 22'h0100011100101100001010;
                12'h07d0: douta_buf <= 22'h1000011100101100001010;
                12'h07d1: douta_buf <= 22'h0100111101001100100010;
                12'h07d2: douta_buf <= 22'h1000111101001100100010;
                12'h07d3: douta_buf <= 22'h0001011101101101000110;
                12'h07d4: douta_buf <= 22'h0101111110001100001010;
                12'h07d5: douta_buf <= 22'h1001111110001100001010;
                12'h07d6: douta_buf <= 22'h0110011110101100100010;
                12'h07d7: douta_buf <= 22'h1010011110101100100010;
                12'h07d8: douta_buf <= 22'h0010111111001101000110;
                12'h07d9: douta_buf <= 22'h0100001100011101000110;
                12'h07da: douta_buf <= 22'h1000001100011101000110;
                12'h07db: douta_buf <= 22'h0100101100111100001010;
                12'h07dc: douta_buf <= 22'h1000101100111100001010;
                12'h07dd: douta_buf <= 22'h0001001101011100100010;
                12'h07de: douta_buf <= 22'h0101101101111101000110;
                12'h07df: douta_buf <= 22'h1001101101111101000110;
                12'h07e0: douta_buf <= 22'h0110001110011100001010;
                12'h07e1: douta_buf <= 22'h1010001110011100001010;
                12'h07e2: douta_buf <= 22'h0010101110111100100010;
                12'h07e3: douta_buf <= 22'h0111001100001101001110;
                12'h07e4: douta_buf <= 22'h1011001100001101001110;
                12'h07e5: douta_buf <= 22'h0100011100101110110010;
                12'h07e6: douta_buf <= 22'h1000011100101110110010;
                12'h07e7: douta_buf <= 22'h0000111101001101110110;
                12'h07e8: douta_buf <= 22'h0101011101101110001110;
                12'h07e9: douta_buf <= 22'h1001011101101110001110;
                12'h07ea: douta_buf <= 22'h0101111110001110110010;
                12'h07eb: douta_buf <= 22'h1001111110001110110010;
                12'h07ec: douta_buf <= 22'h0010011110101101110110;
                12'h07ed: douta_buf <= 22'h0110111111001110001110;
                12'h07ee: douta_buf <= 22'h1010111111001110001110;
                12'h07ef: douta_buf <= 22'h0100001100011110001110;
                12'h07f0: douta_buf <= 22'h1000001100011110001110;
                12'h07f1: douta_buf <= 22'h0000101100111110110010;
                12'h07f2: douta_buf <= 22'h0101001101011101110110;
                12'h07f3: douta_buf <= 22'h1001001101011101110110;
                12'h07f4: douta_buf <= 22'h0101101101111110001110;
                12'h07f5: douta_buf <= 22'h1001101101111110001110;
                12'h07f6: douta_buf <= 22'h0010001110011110110010;
                12'h07f7: douta_buf <= 22'h0110101110111101110110;
                12'h07f8: douta_buf <= 22'h1010101110111101110110;
                12'h07f9: douta_buf <= 22'h0111001100001110010110;
                12'h07fa: douta_buf <= 22'h1011001100001110010110;
                12'h07fb: douta_buf <= 22'h0000011100101110001110;
                12'h07fc: douta_buf <= 22'h0100111101001110110010;
                12'h07fd: douta_buf <= 22'h1000111101001110110010;
                12'h07fe: douta_buf <= 22'h0101011101101101110110;
                12'h07ff: douta_buf <= 22'h1001011101101101110110;
                12'h0800: douta_buf <= 22'h0001111110001110001110;
                12'h0801: douta_buf <= 22'h0110011110101110110010;
                12'h0802: douta_buf <= 22'h1010011110101110110010;
                12'h0803: douta_buf <= 22'h0110111111001101110110;
                12'h0804: douta_buf <= 22'h1010111111001101110110;
                12'h0805: douta_buf <= 22'h0001101000000000000001;
                12'h0806: douta_buf <= 22'h0000000000000000000000;
                12'h0807: douta_buf <= 22'h0000000000000000000000;
                12'h0808: douta_buf <= 22'h0000000000000000000000;
                12'h0809: douta_buf <= 22'h0000000000000000000000;
                12'h080a: douta_buf <= 22'h0000000000000000000000;
                12'h080b: douta_buf <= 22'h0000000000000000000000;
                12'h080c: douta_buf <= 22'h0000000000000000000000;
                12'h080d: douta_buf <= 22'h0000000000000000000000;
                12'h080e: douta_buf <= 22'h0000000000000000000000;
                12'h080f: douta_buf <= 22'h0000000000000000000000;
                12'h0810: douta_buf <= 22'h0000000000000000000000;
                12'h0811: douta_buf <= 22'h0000000000000000000000;
                12'h0812: douta_buf <= 22'h0000000000000000000000;
                12'h0813: douta_buf <= 22'h0000000000000000000000;
                12'h0814: douta_buf <= 22'h0000000000000000000000;
                12'h0815: douta_buf <= 22'h0000000000000000000000;
                12'h0816: douta_buf <= 22'h0000000000000000000000;
                12'h0817: douta_buf <= 22'h0000000000000000000000;
                12'h0818: douta_buf <= 22'h0000000000000000000000;
                12'h0819: douta_buf <= 22'h0000000000000000000000;
                12'h081a: douta_buf <= 22'h0000000000000000000000;
                12'h081b: douta_buf <= 22'h0000000000000000000000;
                12'h081c: douta_buf <= 22'h0000000000000000000000;
                12'h081d: douta_buf <= 22'h0000000000000000000000;
                12'h081e: douta_buf <= 22'h0000000000000000000000;
                12'h081f: douta_buf <= 22'h0000000000000000000000;
                12'h0820: douta_buf <= 22'h0000000000000000000000;
                12'h0821: douta_buf <= 22'h0000000000000000000000;
                12'h0822: douta_buf <= 22'h0000000000000000000000;
                12'h0823: douta_buf <= 22'h0000000000000000000000;
                12'h0824: douta_buf <= 22'h0000000000000000000000;
                12'h0825: douta_buf <= 22'h0000000000000000000000;
                12'h0826: douta_buf <= 22'h0000000000000000000000;
                12'h0827: douta_buf <= 22'h0000000000000000000000;
                12'h0828: douta_buf <= 22'h0000000000000000000000;
                12'h0829: douta_buf <= 22'h0000000000000000000000;
                12'h082a: douta_buf <= 22'h0000000000000000000000;
                12'h082b: douta_buf <= 22'h0000000000000000000000;
                12'h082c: douta_buf <= 22'h0000000000000000000000;
                12'h082d: douta_buf <= 22'h0000000000000000000000;
                12'h082e: douta_buf <= 22'h0000000000000000000000;
                12'h082f: douta_buf <= 22'h0000000000000000000000;
                12'h0830: douta_buf <= 22'h0000000000000000000000;
                12'h0831: douta_buf <= 22'h0000000000000000000000;
                12'h0832: douta_buf <= 22'h0000000000000000000000;
                12'h0833: douta_buf <= 22'h0000000000000000000000;
                12'h0834: douta_buf <= 22'h0000000000000000000000;
                12'h0835: douta_buf <= 22'h0000000000000000000000;
                12'h0836: douta_buf <= 22'h0000000000000000000000;
                12'h0837: douta_buf <= 22'h0000000000000000000000;
                12'h0838: douta_buf <= 22'h0000000000000000000000;
                12'h0839: douta_buf <= 22'h0000000000000000000000;
                12'h083a: douta_buf <= 22'h0000000000000000000000;
                12'h083b: douta_buf <= 22'h0000000000000000000000;
                12'h083c: douta_buf <= 22'h0000000000000000000000;
                12'h083d: douta_buf <= 22'h0000000000000000000000;
                12'h083e: douta_buf <= 22'h0000000000000000000000;
                12'h083f: douta_buf <= 22'h0000000000000000000000;
                12'h0840: douta_buf <= 22'h0000000000000000000000;
                12'h0841: douta_buf <= 22'h0000000000000000000000;
                12'h0842: douta_buf <= 22'h0000000000000000000000;
                12'h0843: douta_buf <= 22'h0000000000000000000000;
                12'h0844: douta_buf <= 22'h0000000000000000000000;
                12'h0845: douta_buf <= 22'h0000000000000000000000;
                12'h0846: douta_buf <= 22'h0000000000000000000000;
                12'h0847: douta_buf <= 22'h0000000000000000000000;
                12'h0848: douta_buf <= 22'h0000000000000000000000;
                12'h0849: douta_buf <= 22'h0000000000000000000000;
                12'h084a: douta_buf <= 22'h0000000000000000000000;
                12'h084b: douta_buf <= 22'h0000000000000000000000;
                12'h084c: douta_buf <= 22'h0000000000000000000000;
                12'h084d: douta_buf <= 22'h0000000000000000000000;
                12'h084e: douta_buf <= 22'h0000000000000000000000;
                12'h084f: douta_buf <= 22'h0000000000000000000000;
                12'h0850: douta_buf <= 22'h0000000000000000000000;
                12'h0851: douta_buf <= 22'h0000000000000000000000;
                12'h0852: douta_buf <= 22'h0000000000000000000000;
                12'h0853: douta_buf <= 22'h0000000000000000000000;
                12'h0854: douta_buf <= 22'h0000000000000000000000;
                12'h0855: douta_buf <= 22'h0000000000000000000000;
                12'h0856: douta_buf <= 22'h0000000000000000000000;
                12'h0857: douta_buf <= 22'h0000000000000000000000;
                12'h0858: douta_buf <= 22'h0000000000000000000000;
                12'h0859: douta_buf <= 22'h0000000000000000000000;
                12'h085a: douta_buf <= 22'h0000000000000000000000;
                12'h085b: douta_buf <= 22'h0000000000000000000000;
                12'h085c: douta_buf <= 22'h0000000000000000000000;
                12'h085d: douta_buf <= 22'h0000000000000000000000;
                12'h085e: douta_buf <= 22'h0000000000000000000000;
                12'h085f: douta_buf <= 22'h0000000000000000000000;
                12'h0860: douta_buf <= 22'h0000000000000000000000;
                12'h0861: douta_buf <= 22'h0000000000000000000000;
                12'h0862: douta_buf <= 22'h0000000000000000000000;
                12'h0863: douta_buf <= 22'h0000000000000000000000;
                12'h0864: douta_buf <= 22'h0000000000000000000000;
                12'h0865: douta_buf <= 22'h0000000000000000000000;
                12'h0866: douta_buf <= 22'h0000000000000000000000;
                12'h0867: douta_buf <= 22'h0000000000000000000000;
                12'h0868: douta_buf <= 22'h0000000000000000000000;
                12'h0869: douta_buf <= 22'h0000000000000000000000;
                12'h086a: douta_buf <= 22'h0000000000000000000000;
                12'h086b: douta_buf <= 22'h0000000000000000000000;
                12'h086c: douta_buf <= 22'h0000000000000000000000;
                12'h086d: douta_buf <= 22'h0000000000000000000000;
                12'h086e: douta_buf <= 22'h0000000000000000000000;
                12'h086f: douta_buf <= 22'h0000000000000000000000;
                12'h0870: douta_buf <= 22'h0000000000000000000000;
                12'h0871: douta_buf <= 22'h0000000000000000000000;
                12'h0872: douta_buf <= 22'h0000000000000000000000;
                12'h0873: douta_buf <= 22'h0000000000000000000000;
                12'h0874: douta_buf <= 22'h0000000000000000000000;
                12'h0875: douta_buf <= 22'h0000000000000000000000;
                12'h0876: douta_buf <= 22'h0000000000000000000000;
                12'h0877: douta_buf <= 22'h0000000000000000000000;
                12'h0878: douta_buf <= 22'h0000000000000000000000;
                12'h0879: douta_buf <= 22'h0000000000000000000000;
                12'h087a: douta_buf <= 22'h0000000000000000000000;
                12'h087b: douta_buf <= 22'h0000000000000000000000;
                12'h087c: douta_buf <= 22'h0000000000000000000000;
                12'h087d: douta_buf <= 22'h0000000000000000000000;
                12'h087e: douta_buf <= 22'h0000000000000000000000;
                12'h087f: douta_buf <= 22'h0000000000000000000000;
                12'h0880: douta_buf <= 22'h0000000000000000000000;
                12'h0881: douta_buf <= 22'h0000000000000000000000;
                12'h0882: douta_buf <= 22'h0000000000000000000000;
                12'h0883: douta_buf <= 22'h0000000000000000000000;
                12'h0884: douta_buf <= 22'h0000000000000000000000;
                12'h0885: douta_buf <= 22'h0000000000000000000000;
                12'h0886: douta_buf <= 22'h0000000000000000000000;
                12'h0887: douta_buf <= 22'h0000000000000000000000;
                12'h0888: douta_buf <= 22'h0000000000000000000000;
                12'h0889: douta_buf <= 22'h0000000000000000000000;
                12'h088a: douta_buf <= 22'h0000000000000000000000;
                12'h088b: douta_buf <= 22'h0000000000000000000000;
                12'h088c: douta_buf <= 22'h0000000000000000000000;
                12'h088d: douta_buf <= 22'h0000000000000000000000;
                12'h088e: douta_buf <= 22'h0000000000000000000000;
                12'h088f: douta_buf <= 22'h0000000000000000000000;
                12'h0890: douta_buf <= 22'h0000000000000000000000;
                12'h0891: douta_buf <= 22'h0000000000000000000000;
                12'h0892: douta_buf <= 22'h0000000000000000000000;
                12'h0893: douta_buf <= 22'h0000000000000000000000;
                12'h0894: douta_buf <= 22'h0000000000000000000000;
                12'h0895: douta_buf <= 22'h0000000000000000000000;
                12'h0896: douta_buf <= 22'h0000000000000000000000;
                12'h0897: douta_buf <= 22'h0000000000000000000000;
                12'h0898: douta_buf <= 22'h0000000000000000000000;
                12'h0899: douta_buf <= 22'h0000000000000000000000;
                12'h089a: douta_buf <= 22'h0000000000000000000000;
                12'h089b: douta_buf <= 22'h0000000000000000000000;
                12'h089c: douta_buf <= 22'h0000000000000000000000;
                12'h089d: douta_buf <= 22'h0000000000000000000000;
                12'h089e: douta_buf <= 22'h0000000000000000000000;
                12'h089f: douta_buf <= 22'h0000000000000000000000;
                12'h08a0: douta_buf <= 22'h0000000000000000000000;
                12'h08a1: douta_buf <= 22'h0000000000000000000000;
                12'h08a2: douta_buf <= 22'h0000000000000000000000;
                12'h08a3: douta_buf <= 22'h0000000000000000000000;
                12'h08a4: douta_buf <= 22'h0000000000000000000000;
                12'h08a5: douta_buf <= 22'h0000000000000000000000;
                12'h08a6: douta_buf <= 22'h0000000000000000000000;
                12'h08a7: douta_buf <= 22'h0000000000000000000000;
                12'h08a8: douta_buf <= 22'h0000000000000000000000;
                12'h08a9: douta_buf <= 22'h0000000000000000000000;
                12'h08aa: douta_buf <= 22'h0000000000000000000000;
                12'h08ab: douta_buf <= 22'h0000000000000000000000;
                12'h08ac: douta_buf <= 22'h0000000000000000000000;
                12'h08ad: douta_buf <= 22'h0000000000000000000000;
                12'h08ae: douta_buf <= 22'h0000000000000000000000;
                12'h08af: douta_buf <= 22'h0000000000000000000000;
                12'h08b0: douta_buf <= 22'h0000000000000000000000;
                12'h08b1: douta_buf <= 22'h0000000000000000000000;
                12'h08b2: douta_buf <= 22'h0000000000000000000000;
                12'h08b3: douta_buf <= 22'h0000000000000000000000;
                12'h08b4: douta_buf <= 22'h0000000000000000000000;
                12'h08b5: douta_buf <= 22'h0000000000000000000000;
                12'h08b6: douta_buf <= 22'h0000000000000000000000;
                12'h08b7: douta_buf <= 22'h0000000000000000000000;
                12'h08b8: douta_buf <= 22'h0000000000000000000000;
                12'h08b9: douta_buf <= 22'h0000000000000000000000;
                12'h08ba: douta_buf <= 22'h0000000000000000000000;
                12'h08bb: douta_buf <= 22'h0000000000000000000000;
                12'h08bc: douta_buf <= 22'h0000000000000000000000;
                12'h08bd: douta_buf <= 22'h0000000000000000000000;
                12'h08be: douta_buf <= 22'h0000000000000000000000;
                12'h08bf: douta_buf <= 22'h0000000000000000000000;
                12'h08c0: douta_buf <= 22'h0000000000000000000000;
                12'h08c1: douta_buf <= 22'h0000000000000000000000;
                12'h08c2: douta_buf <= 22'h0000000000000000000000;
                12'h08c3: douta_buf <= 22'h0000000000000000000000;
                12'h08c4: douta_buf <= 22'h0000000000000000000000;
                12'h08c5: douta_buf <= 22'h0000000000000000000000;
                12'h08c6: douta_buf <= 22'h0000000000000000000000;
                12'h08c7: douta_buf <= 22'h0000000000000000000000;
                12'h08c8: douta_buf <= 22'h0000000000000000000000;
                12'h08c9: douta_buf <= 22'h0000000000000000000000;
                12'h08ca: douta_buf <= 22'h0000000000000000000000;
                12'h08cb: douta_buf <= 22'h0000000000000000000000;
                12'h08cc: douta_buf <= 22'h0000000000000000000000;
                12'h08cd: douta_buf <= 22'h0000000000000000000000;
                12'h08ce: douta_buf <= 22'h0000000000000000000000;
                12'h08cf: douta_buf <= 22'h0000000000000000000000;
                12'h08d0: douta_buf <= 22'h0000000000000000000000;
                12'h08d1: douta_buf <= 22'h0000000000000000000000;
                12'h08d2: douta_buf <= 22'h0000000000000000000000;
                12'h08d3: douta_buf <= 22'h0000000000000000000000;
                12'h08d4: douta_buf <= 22'h0000000000000000000000;
                12'h08d5: douta_buf <= 22'h0000000000000000000000;
                12'h08d6: douta_buf <= 22'h0000000000000000000000;
                12'h08d7: douta_buf <= 22'h0000000000000000000000;
                12'h08d8: douta_buf <= 22'h0000000000000000000000;
                12'h08d9: douta_buf <= 22'h0000000000000000000000;
                12'h08da: douta_buf <= 22'h0000000000000000000000;
                12'h08db: douta_buf <= 22'h0000000000000000000000;
                12'h08dc: douta_buf <= 22'h0000000000000000000000;
                12'h08dd: douta_buf <= 22'h0000000000000000000000;
                12'h08de: douta_buf <= 22'h0000000000000000000000;
                12'h08df: douta_buf <= 22'h0000000000000000000000;
                12'h08e0: douta_buf <= 22'h0000000000000000000000;
                12'h08e1: douta_buf <= 22'h0000000000000000000000;
                12'h08e2: douta_buf <= 22'h0000000000000000000000;
                12'h08e3: douta_buf <= 22'h0000000000000000000000;
                12'h08e4: douta_buf <= 22'h0000000000000000000000;
                12'h08e5: douta_buf <= 22'h0000000000000000000000;
                12'h08e6: douta_buf <= 22'h0000000000000000000000;
                12'h08e7: douta_buf <= 22'h0000000000000000000000;
                12'h08e8: douta_buf <= 22'h0000000000000000000000;
                12'h08e9: douta_buf <= 22'h0000000000000000000000;
                12'h08ea: douta_buf <= 22'h0000000000000000000000;
                12'h08eb: douta_buf <= 22'h0000000000000000000000;
                12'h08ec: douta_buf <= 22'h0000000000000000000000;
                12'h08ed: douta_buf <= 22'h0000000000000000000000;
                12'h08ee: douta_buf <= 22'h0000000000000000000000;
                12'h08ef: douta_buf <= 22'h0000000000000000000000;
                12'h08f0: douta_buf <= 22'h0000000000000000000000;
                12'h08f1: douta_buf <= 22'h0000000000000000000000;
                12'h08f2: douta_buf <= 22'h0000000000000000000000;
                12'h08f3: douta_buf <= 22'h0000000000000000000000;
                12'h08f4: douta_buf <= 22'h0000000000000000000000;
                12'h08f5: douta_buf <= 22'h0000000000000000000000;
                12'h08f6: douta_buf <= 22'h0000000000000000000000;
                12'h08f7: douta_buf <= 22'h0000000000000000000000;
                12'h08f8: douta_buf <= 22'h0000000000000000000000;
                12'h08f9: douta_buf <= 22'h0000000000000000000000;
                12'h08fa: douta_buf <= 22'h0000000000000000000000;
                12'h08fb: douta_buf <= 22'h0000000000000000000000;
                12'h08fc: douta_buf <= 22'h0000000000000000000000;
                12'h08fd: douta_buf <= 22'h0000000000000000000000;
                12'h08fe: douta_buf <= 22'h0000000000000000000000;
                12'h08ff: douta_buf <= 22'h0000000000000000000000;
                12'h0900: douta_buf <= 22'h0000000000000000000000;
                12'h0901: douta_buf <= 22'h0000000000000000000000;
                12'h0902: douta_buf <= 22'h0000000000000000000000;
                12'h0903: douta_buf <= 22'h0000000000000000000000;
                12'h0904: douta_buf <= 22'h0000000000000000000000;
                12'h0905: douta_buf <= 22'h0000000000000000000000;
                12'h0906: douta_buf <= 22'h0000000000000000000000;
                12'h0907: douta_buf <= 22'h0000000000000000000000;
                12'h0908: douta_buf <= 22'h0000000000000000000000;
                12'h0909: douta_buf <= 22'h0000000000000000000000;
                12'h090a: douta_buf <= 22'h0000000000000000000000;
                12'h090b: douta_buf <= 22'h0000000000000000000000;
                12'h090c: douta_buf <= 22'h0000000000000000000000;
                12'h090d: douta_buf <= 22'h0000000000000000000000;
                12'h090e: douta_buf <= 22'h0000000000000000000000;
                12'h090f: douta_buf <= 22'h0000000000000000000000;
                12'h0910: douta_buf <= 22'h0000000000000000000000;
                12'h0911: douta_buf <= 22'h0000000000000000000000;
                12'h0912: douta_buf <= 22'h0000000000000000000000;
                12'h0913: douta_buf <= 22'h0000000000000000000000;
                12'h0914: douta_buf <= 22'h0000000000000000000000;
                12'h0915: douta_buf <= 22'h0000000000000000000000;
                12'h0916: douta_buf <= 22'h0000000000000000000000;
                12'h0917: douta_buf <= 22'h0000000000000000000000;
                12'h0918: douta_buf <= 22'h0000000000000000000000;
                12'h0919: douta_buf <= 22'h0000000000000000000000;
                12'h091a: douta_buf <= 22'h0000000000000000000000;
                12'h091b: douta_buf <= 22'h0000000000000000000000;
                12'h091c: douta_buf <= 22'h0000000000000000000000;
                12'h091d: douta_buf <= 22'h0000000000000000000000;
                12'h091e: douta_buf <= 22'h0000000000000000000000;
                12'h091f: douta_buf <= 22'h0000000000000000000000;
                12'h0920: douta_buf <= 22'h0000000000000000000000;
                12'h0921: douta_buf <= 22'h0000000000000000000000;
                12'h0922: douta_buf <= 22'h0000000000000000000000;
                12'h0923: douta_buf <= 22'h0000000000000000000000;
                12'h0924: douta_buf <= 22'h0000000000000000000000;
                12'h0925: douta_buf <= 22'h0000000000000000000000;
                12'h0926: douta_buf <= 22'h0000000000000000000000;
                12'h0927: douta_buf <= 22'h0000000000000000000000;
                12'h0928: douta_buf <= 22'h0000000000000000000000;
                12'h0929: douta_buf <= 22'h0000000000000000000000;
                12'h092a: douta_buf <= 22'h0000000000000000000000;
                12'h092b: douta_buf <= 22'h0000000000000000000000;
                12'h092c: douta_buf <= 22'h0000000000000000000000;
                12'h092d: douta_buf <= 22'h0000000000000000000000;
                12'h092e: douta_buf <= 22'h0000000000000000000000;
                12'h092f: douta_buf <= 22'h0000000000000000000000;
                12'h0930: douta_buf <= 22'h0000000000000000000000;
                12'h0931: douta_buf <= 22'h0000000000000000000000;
                12'h0932: douta_buf <= 22'h0000000000000000000000;
                12'h0933: douta_buf <= 22'h0000000000000000000000;
                12'h0934: douta_buf <= 22'h0000000000000000000000;
                12'h0935: douta_buf <= 22'h0000000000000000000000;
                12'h0936: douta_buf <= 22'h0000000000000000000000;
                12'h0937: douta_buf <= 22'h0000000000000000000000;
                12'h0938: douta_buf <= 22'h0000000000000000000000;
                12'h0939: douta_buf <= 22'h0000000000000000000000;
                12'h093a: douta_buf <= 22'h0000000000000000000000;
                12'h093b: douta_buf <= 22'h0000000000000000000000;
                12'h093c: douta_buf <= 22'h0000000000000000000000;
                12'h093d: douta_buf <= 22'h0000000000000000000000;
                12'h093e: douta_buf <= 22'h0000000000000000000000;
                12'h093f: douta_buf <= 22'h0000000000000000000000;
                12'h0940: douta_buf <= 22'h0000000000000000000000;
                12'h0941: douta_buf <= 22'h0000000000000000000000;
                12'h0942: douta_buf <= 22'h0000000000000000000000;
                12'h0943: douta_buf <= 22'h0000000000000000000000;
                12'h0944: douta_buf <= 22'h0000000000000000000000;
                12'h0945: douta_buf <= 22'h0000000000000000000000;
                12'h0946: douta_buf <= 22'h0000000000000000000000;
                12'h0947: douta_buf <= 22'h0000000000000000000000;
                12'h0948: douta_buf <= 22'h0000000000000000000000;
                12'h0949: douta_buf <= 22'h0000000000000000000000;
                12'h094a: douta_buf <= 22'h0000000000000000000000;
                12'h094b: douta_buf <= 22'h0000000000000000000000;
                12'h094c: douta_buf <= 22'h0000000000000000000000;
                12'h094d: douta_buf <= 22'h0000000000000000000000;
                12'h094e: douta_buf <= 22'h0000000000000000000000;
                12'h094f: douta_buf <= 22'h0000000000000000000000;
                12'h0950: douta_buf <= 22'h0000000000000000000000;
                12'h0951: douta_buf <= 22'h0000000000000000000000;
                12'h0952: douta_buf <= 22'h0000000000000000000000;
                12'h0953: douta_buf <= 22'h0000000000000000000000;
                12'h0954: douta_buf <= 22'h0000000000000000000000;
                12'h0955: douta_buf <= 22'h0000000000000000000000;
                12'h0956: douta_buf <= 22'h0000000000000000000000;
                12'h0957: douta_buf <= 22'h0000000000000000000000;
                12'h0958: douta_buf <= 22'h0000000000000000000000;
                12'h0959: douta_buf <= 22'h0000000000000000000000;
                12'h095a: douta_buf <= 22'h0000000000000000000000;
                12'h095b: douta_buf <= 22'h0000000000000000000000;
                12'h095c: douta_buf <= 22'h0000000000000000000000;
                12'h095d: douta_buf <= 22'h0000000000000000000000;
                12'h095e: douta_buf <= 22'h0000000000000000000000;
                12'h095f: douta_buf <= 22'h0000000000000000000000;
                12'h0960: douta_buf <= 22'h0000000000000000000000;
                12'h0961: douta_buf <= 22'h0000000000000000000000;
                12'h0962: douta_buf <= 22'h0000000000000000000000;
                12'h0963: douta_buf <= 22'h0000000000000000000000;
                12'h0964: douta_buf <= 22'h0000000000000000000000;
                12'h0965: douta_buf <= 22'h0000000000000000000000;
                12'h0966: douta_buf <= 22'h0000000000000000000000;
                12'h0967: douta_buf <= 22'h0000000000000000000000;
                12'h0968: douta_buf <= 22'h0000000000000000000000;
                12'h0969: douta_buf <= 22'h0000000000000000000000;
                12'h096a: douta_buf <= 22'h0000000000000000000000;
                12'h096b: douta_buf <= 22'h0000000000000000000000;
                12'h096c: douta_buf <= 22'h0000000000000000000000;
                12'h096d: douta_buf <= 22'h0000000000000000000000;
                12'h096e: douta_buf <= 22'h0000000000000000000000;
                12'h096f: douta_buf <= 22'h0000000000000000000000;
                12'h0970: douta_buf <= 22'h0000000000000000000000;
                12'h0971: douta_buf <= 22'h0000000000000000000000;
                12'h0972: douta_buf <= 22'h0000000000000000000000;
                12'h0973: douta_buf <= 22'h0000000000000000000000;
                12'h0974: douta_buf <= 22'h0000000000000000000000;
                12'h0975: douta_buf <= 22'h0000000000000000000000;
                12'h0976: douta_buf <= 22'h0000000000000000000000;
                12'h0977: douta_buf <= 22'h0000000000000000000000;
                12'h0978: douta_buf <= 22'h0000000000000000000000;
                12'h0979: douta_buf <= 22'h0000000000000000000000;
                12'h097a: douta_buf <= 22'h0000000000000000000000;
                12'h097b: douta_buf <= 22'h0000000000000000000000;
                12'h097c: douta_buf <= 22'h0000000000000000000000;
                12'h097d: douta_buf <= 22'h0000000000000000000000;
                12'h097e: douta_buf <= 22'h0000000000000000000000;
                12'h097f: douta_buf <= 22'h0000000000000000000000;
                12'h0980: douta_buf <= 22'h0000000000000000000000;
                12'h0981: douta_buf <= 22'h0000000000000000000000;
                12'h0982: douta_buf <= 22'h0000000000000000000000;
                12'h0983: douta_buf <= 22'h0000000000000000000000;
                12'h0984: douta_buf <= 22'h0000000000000000000000;
                12'h0985: douta_buf <= 22'h0000000000000000000000;
                12'h0986: douta_buf <= 22'h0000000000000000000000;
                12'h0987: douta_buf <= 22'h0000000000000000000000;
                12'h0988: douta_buf <= 22'h0000000000000000000000;
                12'h0989: douta_buf <= 22'h0000000000000000000000;
                12'h098a: douta_buf <= 22'h0000000000000000000000;
                12'h098b: douta_buf <= 22'h0000000000000000000000;
                12'h098c: douta_buf <= 22'h0000000000000000000000;
                12'h098d: douta_buf <= 22'h0000000000000000000000;
                12'h098e: douta_buf <= 22'h0000000000000000000000;
                12'h098f: douta_buf <= 22'h0000000000000000000000;
                12'h0990: douta_buf <= 22'h0000000000000000000000;
                12'h0991: douta_buf <= 22'h0000000000000000000000;
                12'h0992: douta_buf <= 22'h0000000000000000000000;
                12'h0993: douta_buf <= 22'h0000000000000000000000;
                12'h0994: douta_buf <= 22'h0000000000000000000000;
                12'h0995: douta_buf <= 22'h0000000000000000000000;
                12'h0996: douta_buf <= 22'h0000000000000000000000;
                12'h0997: douta_buf <= 22'h0000000000000000000000;
                12'h0998: douta_buf <= 22'h0000000000000000000000;
                12'h0999: douta_buf <= 22'h0000000000000000000000;
                12'h099a: douta_buf <= 22'h0000000000000000000000;
                12'h099b: douta_buf <= 22'h0000000000000000000000;
                12'h099c: douta_buf <= 22'h0000000000000000000000;
                12'h099d: douta_buf <= 22'h0000000000000000000000;
                12'h099e: douta_buf <= 22'h0000000000000000000000;
                12'h099f: douta_buf <= 22'h0000000000000000000000;
                12'h09a0: douta_buf <= 22'h0000000000000000000000;
                12'h09a1: douta_buf <= 22'h0000000000000000000000;
                12'h09a2: douta_buf <= 22'h0000000000000000000000;
                12'h09a3: douta_buf <= 22'h0000000000000000000000;
                12'h09a4: douta_buf <= 22'h0000000000000000000000;
                12'h09a5: douta_buf <= 22'h0000000000000000000000;
                12'h09a6: douta_buf <= 22'h0000000000000000000000;
                12'h09a7: douta_buf <= 22'h0000000000000000000000;
                12'h09a8: douta_buf <= 22'h0000000000000000000000;
                12'h09a9: douta_buf <= 22'h0000000000000000000000;
                12'h09aa: douta_buf <= 22'h0000000000000000000000;
                12'h09ab: douta_buf <= 22'h0000000000000000000000;
                12'h09ac: douta_buf <= 22'h0000000000000000000000;
                12'h09ad: douta_buf <= 22'h0000000000000000000000;
                12'h09ae: douta_buf <= 22'h0000000000000000000000;
                12'h09af: douta_buf <= 22'h0000000000000000000000;
                12'h09b0: douta_buf <= 22'h0000000000000000000000;
                12'h09b1: douta_buf <= 22'h0000000000000000000000;
                12'h09b2: douta_buf <= 22'h0000000000000000000000;
                12'h09b3: douta_buf <= 22'h0000000000000000000000;
                12'h09b4: douta_buf <= 22'h0000000000000000000000;
                12'h09b5: douta_buf <= 22'h0000000000000000000000;
                12'h09b6: douta_buf <= 22'h0000000000000000000000;
                12'h09b7: douta_buf <= 22'h0000000000000000000000;
                12'h09b8: douta_buf <= 22'h0000000000000000000000;
                12'h09b9: douta_buf <= 22'h0000000000000000000000;
                12'h09ba: douta_buf <= 22'h0000000000000000000000;
                12'h09bb: douta_buf <= 22'h0000000000000000000000;
                12'h09bc: douta_buf <= 22'h0000000000000000000000;
                12'h09bd: douta_buf <= 22'h0000000000000000000000;
                12'h09be: douta_buf <= 22'h0000000000000000000000;
                12'h09bf: douta_buf <= 22'h0000000000000000000000;
                12'h09c0: douta_buf <= 22'h0000000000000000000000;
                12'h09c1: douta_buf <= 22'h0000000000000000000000;
                12'h09c2: douta_buf <= 22'h0000000000000000000000;
                12'h09c3: douta_buf <= 22'h0000000000000000000000;
                12'h09c4: douta_buf <= 22'h0000000000000000000000;
                12'h09c5: douta_buf <= 22'h0000000000000000000000;
                12'h09c6: douta_buf <= 22'h0000000000000000000000;
                12'h09c7: douta_buf <= 22'h0000000000000000000000;
                12'h09c8: douta_buf <= 22'h0000000000000000000000;
                12'h09c9: douta_buf <= 22'h0000000000000000000000;
                12'h09ca: douta_buf <= 22'h0000000000000000000000;
                12'h09cb: douta_buf <= 22'h0000000000000000000000;
                12'h09cc: douta_buf <= 22'h0000000000000000000000;
                12'h09cd: douta_buf <= 22'h0000000000000000000000;
                12'h09ce: douta_buf <= 22'h0000000000000000000000;
                12'h09cf: douta_buf <= 22'h0000000000000000000000;
                12'h09d0: douta_buf <= 22'h0000000000000000000000;
                12'h09d1: douta_buf <= 22'h0000000000000000000000;
                12'h09d2: douta_buf <= 22'h0000000000000000000000;
                12'h09d3: douta_buf <= 22'h0000000000000000000000;
                12'h09d4: douta_buf <= 22'h0000000000000000000000;
                12'h09d5: douta_buf <= 22'h0000000000000000000000;
                12'h09d6: douta_buf <= 22'h0000000000000000000000;
                12'h09d7: douta_buf <= 22'h0000000000000000000000;
                12'h09d8: douta_buf <= 22'h0000000000000000000000;
                12'h09d9: douta_buf <= 22'h0000000000000000000000;
                12'h09da: douta_buf <= 22'h0000000000000000000000;
                12'h09db: douta_buf <= 22'h0000000000000000000000;
                12'h09dc: douta_buf <= 22'h0000000000000000000000;
                12'h09dd: douta_buf <= 22'h0000000000000000000000;
                12'h09de: douta_buf <= 22'h0000000000000000000000;
                12'h09df: douta_buf <= 22'h0000000000000000000000;
                12'h09e0: douta_buf <= 22'h0000000000000000000000;
                12'h09e1: douta_buf <= 22'h0000000000000000000000;
                12'h09e2: douta_buf <= 22'h0000000000000000000000;
                12'h09e3: douta_buf <= 22'h0000000000000000000000;
                12'h09e4: douta_buf <= 22'h0000000000000000000000;
                12'h09e5: douta_buf <= 22'h0000000000000000000000;
                12'h09e6: douta_buf <= 22'h0000000000000000000000;
                12'h09e7: douta_buf <= 22'h0000000000000000000000;
                12'h09e8: douta_buf <= 22'h0000000000000000000000;
                12'h09e9: douta_buf <= 22'h0000000000000000000000;
                12'h09ea: douta_buf <= 22'h0000000000000000000000;
                12'h09eb: douta_buf <= 22'h0000000000000000000000;
                12'h09ec: douta_buf <= 22'h0000000000000000000000;
                12'h09ed: douta_buf <= 22'h0000000000000000000000;
                12'h09ee: douta_buf <= 22'h0000000000000000000000;
                12'h09ef: douta_buf <= 22'h0000000000000000000000;
                12'h09f0: douta_buf <= 22'h0000000000000000000000;
                12'h09f1: douta_buf <= 22'h0000000000000000000000;
                12'h09f2: douta_buf <= 22'h0000000000000000000000;
                12'h09f3: douta_buf <= 22'h0000000000000000000000;
                12'h09f4: douta_buf <= 22'h0000000000000000000000;
                12'h09f5: douta_buf <= 22'h0000000000000000000000;
                12'h09f6: douta_buf <= 22'h0000000000000000000000;
                12'h09f7: douta_buf <= 22'h0000000000000000000000;
                12'h09f8: douta_buf <= 22'h0000000000000000000000;
                12'h09f9: douta_buf <= 22'h0000000000000000000000;
                12'h09fa: douta_buf <= 22'h0000000000000000000000;
                12'h09fb: douta_buf <= 22'h0000000000000000000000;
                12'h09fc: douta_buf <= 22'h0000000000000000000000;
                12'h09fd: douta_buf <= 22'h0000000000000000000000;
                12'h09fe: douta_buf <= 22'h0000000000000000000000;
                12'h09ff: douta_buf <= 22'h0000000000000000000000;
                12'h0a00: douta_buf <= 22'h0000000000000000000000;
                12'h0a01: douta_buf <= 22'h0000000000000000000000;
                12'h0a02: douta_buf <= 22'h0000000000000000000000;
                12'h0a03: douta_buf <= 22'h0000000000000000000000;
                12'h0a04: douta_buf <= 22'h0000000000000000000000;
                12'h0a05: douta_buf <= 22'h0000000000000000000000;
                12'h0a06: douta_buf <= 22'h0000000000000000000000;
                12'h0a07: douta_buf <= 22'h0000000000000000000000;
                12'h0a08: douta_buf <= 22'h0000000000000000000000;
                12'h0a09: douta_buf <= 22'h0000000000000000000000;
                12'h0a0a: douta_buf <= 22'h0000000000000000000000;
                12'h0a0b: douta_buf <= 22'h0000000000000000000000;
                12'h0a0c: douta_buf <= 22'h0000000000000000000000;
                12'h0a0d: douta_buf <= 22'h0000000000000000000000;
                12'h0a0e: douta_buf <= 22'h0000000000000000000000;
                12'h0a0f: douta_buf <= 22'h0000000000000000000000;
                12'h0a10: douta_buf <= 22'h0000000000000000000000;
                12'h0a11: douta_buf <= 22'h0000000000000000000000;
                12'h0a12: douta_buf <= 22'h0000000000000000000000;
                12'h0a13: douta_buf <= 22'h0000000000000000000000;
                12'h0a14: douta_buf <= 22'h0000000000000000000000;
                12'h0a15: douta_buf <= 22'h0000000000000000000000;
                12'h0a16: douta_buf <= 22'h0000000000000000000000;
                12'h0a17: douta_buf <= 22'h0000000000000000000000;
                12'h0a18: douta_buf <= 22'h0000000000000000000000;
                12'h0a19: douta_buf <= 22'h0000000000000000000000;
                12'h0a1a: douta_buf <= 22'h0000000000000000000000;
                12'h0a1b: douta_buf <= 22'h0000000000000000000000;
                12'h0a1c: douta_buf <= 22'h0000000000000000000000;
                12'h0a1d: douta_buf <= 22'h0000000000000000000000;
                12'h0a1e: douta_buf <= 22'h0000000000000000000000;
                12'h0a1f: douta_buf <= 22'h0000000000000000000000;
                12'h0a20: douta_buf <= 22'h0000000000000000000000;
                12'h0a21: douta_buf <= 22'h0000000000000000000000;
                12'h0a22: douta_buf <= 22'h0000000000000000000000;
                12'h0a23: douta_buf <= 22'h0000000000000000000000;
                12'h0a24: douta_buf <= 22'h0000000000000000000000;
                12'h0a25: douta_buf <= 22'h0000000000000000000000;
                12'h0a26: douta_buf <= 22'h0000000000000000000000;
                12'h0a27: douta_buf <= 22'h0000000000000000000000;
                12'h0a28: douta_buf <= 22'h0000000000000000000000;
                12'h0a29: douta_buf <= 22'h0000000000000000000000;
                12'h0a2a: douta_buf <= 22'h0000000000000000000000;
                12'h0a2b: douta_buf <= 22'h0000000000000000000000;
                12'h0a2c: douta_buf <= 22'h0000000000000000000000;
                12'h0a2d: douta_buf <= 22'h0000000000000000000000;
                12'h0a2e: douta_buf <= 22'h0000000000000000000000;
                12'h0a2f: douta_buf <= 22'h0000000000000000000000;
                12'h0a30: douta_buf <= 22'h0000000000000000000000;
                12'h0a31: douta_buf <= 22'h0000000000000000000000;
                12'h0a32: douta_buf <= 22'h0000000000000000000000;
                12'h0a33: douta_buf <= 22'h0000000000000000000000;
                12'h0a34: douta_buf <= 22'h0000000000000000000000;
                12'h0a35: douta_buf <= 22'h0000000000000000000000;
                12'h0a36: douta_buf <= 22'h0000000000000000000000;
                12'h0a37: douta_buf <= 22'h0000000000000000000000;
                12'h0a38: douta_buf <= 22'h0000000000000000000000;
                12'h0a39: douta_buf <= 22'h0000000000000000000000;
                12'h0a3a: douta_buf <= 22'h0000000000000000000000;
                12'h0a3b: douta_buf <= 22'h0000000000000000000000;
                12'h0a3c: douta_buf <= 22'h0000000000000000000000;
                12'h0a3d: douta_buf <= 22'h0000000000000000000000;
                12'h0a3e: douta_buf <= 22'h0000000000000000000000;
                12'h0a3f: douta_buf <= 22'h0000000000000000000000;
                12'h0a40: douta_buf <= 22'h0000000000000000000000;
                12'h0a41: douta_buf <= 22'h0000000000000000000000;
                12'h0a42: douta_buf <= 22'h0000000000000000000000;
                12'h0a43: douta_buf <= 22'h0000000000000000000000;
                12'h0a44: douta_buf <= 22'h0000000000000000000000;
                12'h0a45: douta_buf <= 22'h0000000000000000000000;
                12'h0a46: douta_buf <= 22'h0000000000000000000000;
                12'h0a47: douta_buf <= 22'h0000000000000000000000;
                12'h0a48: douta_buf <= 22'h0000000000000000000000;
                12'h0a49: douta_buf <= 22'h0000000000000000000000;
                12'h0a4a: douta_buf <= 22'h0000000000000000000000;
                12'h0a4b: douta_buf <= 22'h0000000000000000000000;
                12'h0a4c: douta_buf <= 22'h0000000000000000000000;
                12'h0a4d: douta_buf <= 22'h0000000000000000000000;
                12'h0a4e: douta_buf <= 22'h0000000000000000000000;
                12'h0a4f: douta_buf <= 22'h0000000000000000000000;
                12'h0a50: douta_buf <= 22'h0000000000000000000000;
                12'h0a51: douta_buf <= 22'h0000000000000000000000;
                12'h0a52: douta_buf <= 22'h0000000000000000000000;
                12'h0a53: douta_buf <= 22'h0000000000000000000000;
                12'h0a54: douta_buf <= 22'h0000000000000000000000;
                12'h0a55: douta_buf <= 22'h0000000000000000000000;
                12'h0a56: douta_buf <= 22'h0000000000000000000000;
                12'h0a57: douta_buf <= 22'h0000000000000000000000;
                12'h0a58: douta_buf <= 22'h0000000000000000000000;
                12'h0a59: douta_buf <= 22'h0000000000000000000000;
                12'h0a5a: douta_buf <= 22'h0000000000000000000000;
                12'h0a5b: douta_buf <= 22'h0000000000000000000000;
                12'h0a5c: douta_buf <= 22'h0000000000000000000000;
                12'h0a5d: douta_buf <= 22'h0000000000000000000000;
                12'h0a5e: douta_buf <= 22'h0000000000000000000000;
                12'h0a5f: douta_buf <= 22'h0000000000000000000000;
                12'h0a60: douta_buf <= 22'h0000000000000000000000;
                12'h0a61: douta_buf <= 22'h0000000000000000000000;
                12'h0a62: douta_buf <= 22'h0000000000000000000000;
                12'h0a63: douta_buf <= 22'h0000000000000000000000;
                12'h0a64: douta_buf <= 22'h0000000000000000000000;
                12'h0a65: douta_buf <= 22'h0000000000000000000000;
                12'h0a66: douta_buf <= 22'h0000000000000000000000;
                12'h0a67: douta_buf <= 22'h0000000000000000000000;
                12'h0a68: douta_buf <= 22'h0000000000000000000000;
                12'h0a69: douta_buf <= 22'h0000000000000000000000;
                12'h0a6a: douta_buf <= 22'h0000000000000000000000;
                12'h0a6b: douta_buf <= 22'h0000000000000000000000;
                12'h0a6c: douta_buf <= 22'h0000000000000000000000;
                12'h0a6d: douta_buf <= 22'h0000000000000000000000;
                12'h0a6e: douta_buf <= 22'h0000000000000000000000;
                12'h0a6f: douta_buf <= 22'h0000000000000000000000;
                12'h0a70: douta_buf <= 22'h0000000000000000000000;
                12'h0a71: douta_buf <= 22'h0000000000000000000000;
                12'h0a72: douta_buf <= 22'h0000000000000000000000;
                12'h0a73: douta_buf <= 22'h0000000000000000000000;
                12'h0a74: douta_buf <= 22'h0000000000000000000000;
                12'h0a75: douta_buf <= 22'h0000000000000000000000;
                12'h0a76: douta_buf <= 22'h0000000000000000000000;
                12'h0a77: douta_buf <= 22'h0000000000000000000000;
                12'h0a78: douta_buf <= 22'h0000000000000000000000;
                12'h0a79: douta_buf <= 22'h0000000000000000000000;
                12'h0a7a: douta_buf <= 22'h0000000000000000000000;
                12'h0a7b: douta_buf <= 22'h0000000000000000000000;
                12'h0a7c: douta_buf <= 22'h0000000000000000000000;
                12'h0a7d: douta_buf <= 22'h0000000000000000000000;
                12'h0a7e: douta_buf <= 22'h0000000000000000000000;
                12'h0a7f: douta_buf <= 22'h0000000000000000000000;
                12'h0a80: douta_buf <= 22'h0000000000000000000000;
                12'h0a81: douta_buf <= 22'h0000000000000000000000;
                12'h0a82: douta_buf <= 22'h0000000000000000000000;
                12'h0a83: douta_buf <= 22'h0000000000000000000000;
                12'h0a84: douta_buf <= 22'h0000000000000000000000;
                12'h0a85: douta_buf <= 22'h0000000000000000000000;
                12'h0a86: douta_buf <= 22'h0000000000000000000000;
                12'h0a87: douta_buf <= 22'h0000000000000000000000;
                12'h0a88: douta_buf <= 22'h0000000000000000000000;
                12'h0a89: douta_buf <= 22'h0000000000000000000000;
                12'h0a8a: douta_buf <= 22'h0000000000000000000000;
                12'h0a8b: douta_buf <= 22'h0000000000000000000000;
                12'h0a8c: douta_buf <= 22'h0000000000000000000000;
                12'h0a8d: douta_buf <= 22'h0000000000000000000000;
                12'h0a8e: douta_buf <= 22'h0000000000000000000000;
                12'h0a8f: douta_buf <= 22'h0000000000000000000000;
                12'h0a90: douta_buf <= 22'h0000000000000000000000;
                12'h0a91: douta_buf <= 22'h0000000000000000000000;
                12'h0a92: douta_buf <= 22'h0000000000000000000000;
                12'h0a93: douta_buf <= 22'h0000000000000000000000;
                12'h0a94: douta_buf <= 22'h0000000000000000000000;
                12'h0a95: douta_buf <= 22'h0000000000000000000000;
                12'h0a96: douta_buf <= 22'h0000000000000000000000;
                12'h0a97: douta_buf <= 22'h0000000000000000000000;
                12'h0a98: douta_buf <= 22'h0000000000000000000000;
                12'h0a99: douta_buf <= 22'h0000000000000000000000;
                12'h0a9a: douta_buf <= 22'h0000000000000000000000;
                12'h0a9b: douta_buf <= 22'h0000000000000000000000;
                12'h0a9c: douta_buf <= 22'h0000000000000000000000;
                12'h0a9d: douta_buf <= 22'h0000000000000000000000;
                12'h0a9e: douta_buf <= 22'h0000000000000000000000;
                12'h0a9f: douta_buf <= 22'h0000000000000000000000;
                12'h0aa0: douta_buf <= 22'h0000000000000000000000;
                12'h0aa1: douta_buf <= 22'h0000000000000000000000;
                12'h0aa2: douta_buf <= 22'h0000000000000000000000;
                12'h0aa3: douta_buf <= 22'h0000000000000000000000;
                12'h0aa4: douta_buf <= 22'h0000000000000000000000;
                12'h0aa5: douta_buf <= 22'h0000000000000000000000;
                12'h0aa6: douta_buf <= 22'h0000000000000000000000;
                12'h0aa7: douta_buf <= 22'h0000000000000000000000;
                12'h0aa8: douta_buf <= 22'h0000000000000000000000;
                12'h0aa9: douta_buf <= 22'h0000000000000000000000;
                12'h0aaa: douta_buf <= 22'h0000000000000000000000;
                12'h0aab: douta_buf <= 22'h0000000000000000000000;
                12'h0aac: douta_buf <= 22'h0000000000000000000000;
                12'h0aad: douta_buf <= 22'h0000000000000000000000;
                12'h0aae: douta_buf <= 22'h0000000000000000000000;
                12'h0aaf: douta_buf <= 22'h0000000000000000000000;
                12'h0ab0: douta_buf <= 22'h0000000000000000000000;
                12'h0ab1: douta_buf <= 22'h0000000000000000000000;
                12'h0ab2: douta_buf <= 22'h0000000000000000000000;
                12'h0ab3: douta_buf <= 22'h0000000000000000000000;
                12'h0ab4: douta_buf <= 22'h0000000000000000000000;
                12'h0ab5: douta_buf <= 22'h0000000000000000000000;
                12'h0ab6: douta_buf <= 22'h0000000000000000000000;
                12'h0ab7: douta_buf <= 22'h0000000000000000000000;
                12'h0ab8: douta_buf <= 22'h0000000000000000000000;
                12'h0ab9: douta_buf <= 22'h0000000000000000000000;
                12'h0aba: douta_buf <= 22'h0000000000000000000000;
                12'h0abb: douta_buf <= 22'h0000000000000000000000;
                12'h0abc: douta_buf <= 22'h0000000000000000000000;
                12'h0abd: douta_buf <= 22'h0000000000000000000000;
                12'h0abe: douta_buf <= 22'h0000000000000000000000;
                12'h0abf: douta_buf <= 22'h0000000000000000000000;
                12'h0ac0: douta_buf <= 22'h0000000000000000000000;
                12'h0ac1: douta_buf <= 22'h0000000000000000000000;
                12'h0ac2: douta_buf <= 22'h0000000000000000000000;
                12'h0ac3: douta_buf <= 22'h0000000000000000000000;
                12'h0ac4: douta_buf <= 22'h0000000000000000000000;
                12'h0ac5: douta_buf <= 22'h0000000000000000000000;
                12'h0ac6: douta_buf <= 22'h0000000000000000000000;
                12'h0ac7: douta_buf <= 22'h0000000000000000000000;
                12'h0ac8: douta_buf <= 22'h0000000000000000000000;
                12'h0ac9: douta_buf <= 22'h0000000000000000000000;
                12'h0aca: douta_buf <= 22'h0000000000000000000000;
                12'h0acb: douta_buf <= 22'h0000000000000000000000;
                12'h0acc: douta_buf <= 22'h0000000000000000000000;
                12'h0acd: douta_buf <= 22'h0000000000000000000000;
                12'h0ace: douta_buf <= 22'h0000000000000000000000;
                12'h0acf: douta_buf <= 22'h0000000000000000000000;
                12'h0ad0: douta_buf <= 22'h0000000000000000000000;
                12'h0ad1: douta_buf <= 22'h0000000000000000000000;
                12'h0ad2: douta_buf <= 22'h0000000000000000000000;
                12'h0ad3: douta_buf <= 22'h0000000000000000000000;
                12'h0ad4: douta_buf <= 22'h0000000000000000000000;
                12'h0ad5: douta_buf <= 22'h0000000000000000000000;
                12'h0ad6: douta_buf <= 22'h0000000000000000000000;
                12'h0ad7: douta_buf <= 22'h0000000000000000000000;
                12'h0ad8: douta_buf <= 22'h0000000000000000000000;
                12'h0ad9: douta_buf <= 22'h0000000000000000000000;
                12'h0ada: douta_buf <= 22'h0000000000000000000000;
                12'h0adb: douta_buf <= 22'h0000000000000000000000;
                12'h0adc: douta_buf <= 22'h0000000000000000000000;
                12'h0add: douta_buf <= 22'h0000000000000000000000;
                12'h0ade: douta_buf <= 22'h0000000000000000000000;
                12'h0adf: douta_buf <= 22'h0000000000000000000000;
                12'h0ae0: douta_buf <= 22'h0000000000000000000000;
                12'h0ae1: douta_buf <= 22'h0000000000000000000000;
                12'h0ae2: douta_buf <= 22'h0000000000000000000000;
                12'h0ae3: douta_buf <= 22'h0000000000000000000000;
                12'h0ae4: douta_buf <= 22'h0000000000000000000000;
                12'h0ae5: douta_buf <= 22'h0000000000000000000000;
                12'h0ae6: douta_buf <= 22'h0000000000000000000000;
                12'h0ae7: douta_buf <= 22'h0000000000000000000000;
                12'h0ae8: douta_buf <= 22'h0000000000000000000000;
                12'h0ae9: douta_buf <= 22'h0000000000000000000000;
                12'h0aea: douta_buf <= 22'h0000000000000000000000;
                12'h0aeb: douta_buf <= 22'h0000000000000000000000;
                12'h0aec: douta_buf <= 22'h0000000000000000000000;
                12'h0aed: douta_buf <= 22'h0000000000000000000000;
                12'h0aee: douta_buf <= 22'h0000000000000000000000;
                12'h0aef: douta_buf <= 22'h0000000000000000000000;
                12'h0af0: douta_buf <= 22'h0000000000000000000000;
                12'h0af1: douta_buf <= 22'h0000000000000000000000;
                12'h0af2: douta_buf <= 22'h0000000000000000000000;
                12'h0af3: douta_buf <= 22'h0000000000000000000000;
                12'h0af4: douta_buf <= 22'h0000000000000000000000;
                12'h0af5: douta_buf <= 22'h0000000000000000000000;
                12'h0af6: douta_buf <= 22'h0000000000000000000000;
                12'h0af7: douta_buf <= 22'h0000000000000000000000;
                12'h0af8: douta_buf <= 22'h0000000000000000000000;
                12'h0af9: douta_buf <= 22'h0000000000000000000000;
                12'h0afa: douta_buf <= 22'h0000000000000000000000;
                12'h0afb: douta_buf <= 22'h0000000000000000000000;
                12'h0afc: douta_buf <= 22'h0000000000000000000000;
                12'h0afd: douta_buf <= 22'h0000000000000000000000;
                12'h0afe: douta_buf <= 22'h0000000000000000000000;
                12'h0aff: douta_buf <= 22'h0000000000000000000000;
                12'h0b00: douta_buf <= 22'h0000000000000000000000;
                12'h0b01: douta_buf <= 22'h0000000000000000000000;
                12'h0b02: douta_buf <= 22'h0000000000000000000000;
                12'h0b03: douta_buf <= 22'h0000000000000000000000;
                12'h0b04: douta_buf <= 22'h0000000000000000000000;
                12'h0b05: douta_buf <= 22'h0000000000000000000000;
                12'h0b06: douta_buf <= 22'h0000000000000000000000;
                12'h0b07: douta_buf <= 22'h0000000000000000000000;
                12'h0b08: douta_buf <= 22'h0000000000000000000000;
                12'h0b09: douta_buf <= 22'h0000000000000000000000;
                12'h0b0a: douta_buf <= 22'h0000000000000000000000;
                12'h0b0b: douta_buf <= 22'h0000000000000000000000;
                12'h0b0c: douta_buf <= 22'h0000000000000000000000;
                12'h0b0d: douta_buf <= 22'h0000000000000000000000;
                12'h0b0e: douta_buf <= 22'h0000000000000000000000;
                12'h0b0f: douta_buf <= 22'h0000000000000000000000;
                12'h0b10: douta_buf <= 22'h0000000000000000000000;
                12'h0b11: douta_buf <= 22'h0000000000000000000000;
                12'h0b12: douta_buf <= 22'h0000000000000000000000;
                12'h0b13: douta_buf <= 22'h0000000000000000000000;
                12'h0b14: douta_buf <= 22'h0000000000000000000000;
                12'h0b15: douta_buf <= 22'h0000000000000000000000;
                12'h0b16: douta_buf <= 22'h0000000000000000000000;
                12'h0b17: douta_buf <= 22'h0000000000000000000000;
                12'h0b18: douta_buf <= 22'h0000000000000000000000;
                12'h0b19: douta_buf <= 22'h0000000000000000000000;
                12'h0b1a: douta_buf <= 22'h0000000000000000000000;
                12'h0b1b: douta_buf <= 22'h0000000000000000000000;
                12'h0b1c: douta_buf <= 22'h0000000000000000000000;
                12'h0b1d: douta_buf <= 22'h0000000000000000000000;
                12'h0b1e: douta_buf <= 22'h0000000000000000000000;
                12'h0b1f: douta_buf <= 22'h0000000000000000000000;
                12'h0b20: douta_buf <= 22'h0000000000000000000000;
                12'h0b21: douta_buf <= 22'h0000000000000000000000;
                12'h0b22: douta_buf <= 22'h0000000000000000000000;
                12'h0b23: douta_buf <= 22'h0000000000000000000000;
                12'h0b24: douta_buf <= 22'h0000000000000000000000;
                12'h0b25: douta_buf <= 22'h0000000000000000000000;
                12'h0b26: douta_buf <= 22'h0000000000000000000000;
                12'h0b27: douta_buf <= 22'h0000000000000000000000;
                12'h0b28: douta_buf <= 22'h0000000000000000000000;
                12'h0b29: douta_buf <= 22'h0000000000000000000000;
                12'h0b2a: douta_buf <= 22'h0000000000000000000000;
                12'h0b2b: douta_buf <= 22'h0000000000000000000000;
                12'h0b2c: douta_buf <= 22'h0000000000000000000000;
                12'h0b2d: douta_buf <= 22'h0000000000000000000000;
                12'h0b2e: douta_buf <= 22'h0000000000000000000000;
                12'h0b2f: douta_buf <= 22'h0000000000000000000000;
                12'h0b30: douta_buf <= 22'h0000000000000000000000;
                12'h0b31: douta_buf <= 22'h0000000000000000000000;
                12'h0b32: douta_buf <= 22'h0000000000000000000000;
                12'h0b33: douta_buf <= 22'h0000000000000000000000;
                12'h0b34: douta_buf <= 22'h0000000000000000000000;
                12'h0b35: douta_buf <= 22'h0000000000000000000000;
                12'h0b36: douta_buf <= 22'h0000000000000000000000;
                12'h0b37: douta_buf <= 22'h0000000000000000000000;
                12'h0b38: douta_buf <= 22'h0000000000000000000000;
                12'h0b39: douta_buf <= 22'h0000000000000000000000;
                12'h0b3a: douta_buf <= 22'h0000000000000000000000;
                12'h0b3b: douta_buf <= 22'h0000000000000000000000;
                12'h0b3c: douta_buf <= 22'h0000000000000000000000;
                12'h0b3d: douta_buf <= 22'h0000000000000000000000;
                12'h0b3e: douta_buf <= 22'h0000000000000000000000;
                12'h0b3f: douta_buf <= 22'h0000000000000000000000;
                12'h0b40: douta_buf <= 22'h0000000000000000000000;
                12'h0b41: douta_buf <= 22'h0000000000000000000000;
                12'h0b42: douta_buf <= 22'h0000000000000000000000;
                12'h0b43: douta_buf <= 22'h0000000000000000000000;
                12'h0b44: douta_buf <= 22'h0000000000000000000000;
                12'h0b45: douta_buf <= 22'h0000000000000000000000;
                12'h0b46: douta_buf <= 22'h0000000000000000000000;
                12'h0b47: douta_buf <= 22'h0000000000000000000000;
                12'h0b48: douta_buf <= 22'h0000000000000000000000;
                12'h0b49: douta_buf <= 22'h0000000000000000000000;
                12'h0b4a: douta_buf <= 22'h0000000000000000000000;
                12'h0b4b: douta_buf <= 22'h0000000000000000000000;
                12'h0b4c: douta_buf <= 22'h0000000000000000000000;
                12'h0b4d: douta_buf <= 22'h0000000000000000000000;
                12'h0b4e: douta_buf <= 22'h0000000000000000000000;
                12'h0b4f: douta_buf <= 22'h0000000000000000000000;
                12'h0b50: douta_buf <= 22'h0000000000000000000000;
                12'h0b51: douta_buf <= 22'h0000000000000000000000;
                12'h0b52: douta_buf <= 22'h0000000000000000000000;
                12'h0b53: douta_buf <= 22'h0000000000000000000000;
                12'h0b54: douta_buf <= 22'h0000000000000000000000;
                12'h0b55: douta_buf <= 22'h0000000000000000000000;
                12'h0b56: douta_buf <= 22'h0000000000000000000000;
                12'h0b57: douta_buf <= 22'h0000000000000000000000;
                12'h0b58: douta_buf <= 22'h0000000000000000000000;
                12'h0b59: douta_buf <= 22'h0000000000000000000000;
                12'h0b5a: douta_buf <= 22'h0000000000000000000000;
                12'h0b5b: douta_buf <= 22'h0000000000000000000000;
                12'h0b5c: douta_buf <= 22'h0000000000000000000000;
                12'h0b5d: douta_buf <= 22'h0000000000000000000000;
                12'h0b5e: douta_buf <= 22'h0000000000000000000000;
                12'h0b5f: douta_buf <= 22'h0000000000000000000000;
                12'h0b60: douta_buf <= 22'h0000000000000000000000;
                12'h0b61: douta_buf <= 22'h0000000000000000000000;
                12'h0b62: douta_buf <= 22'h0000000000000000000000;
                12'h0b63: douta_buf <= 22'h0000000000000000000000;
                12'h0b64: douta_buf <= 22'h0000000000000000000000;
                12'h0b65: douta_buf <= 22'h0000000000000000000000;
                12'h0b66: douta_buf <= 22'h0000000000000000000000;
                12'h0b67: douta_buf <= 22'h0000000000000000000000;
                12'h0b68: douta_buf <= 22'h0000000000000000000000;
                12'h0b69: douta_buf <= 22'h0000000000000000000000;
                12'h0b6a: douta_buf <= 22'h0000000000000000000000;
                12'h0b6b: douta_buf <= 22'h0000000000000000000000;
                12'h0b6c: douta_buf <= 22'h0000000000000000000000;
                12'h0b6d: douta_buf <= 22'h0000000000000000000000;
                12'h0b6e: douta_buf <= 22'h0000000000000000000000;
                12'h0b6f: douta_buf <= 22'h0000000000000000000000;
                12'h0b70: douta_buf <= 22'h0000000000000000000000;
                12'h0b71: douta_buf <= 22'h0000000000000000000000;
                12'h0b72: douta_buf <= 22'h0000000000000000000000;
                12'h0b73: douta_buf <= 22'h0000000000000000000000;
                12'h0b74: douta_buf <= 22'h0000000000000000000000;
                12'h0b75: douta_buf <= 22'h0000000000000000000000;
                12'h0b76: douta_buf <= 22'h0000000000000000000000;
                12'h0b77: douta_buf <= 22'h0000000000000000000000;
                12'h0b78: douta_buf <= 22'h0000000000000000000000;
                12'h0b79: douta_buf <= 22'h0000000000000000000000;
                12'h0b7a: douta_buf <= 22'h0000000000000000000000;
                12'h0b7b: douta_buf <= 22'h0000000000000000000000;
                12'h0b7c: douta_buf <= 22'h0000000000000000000000;
                12'h0b7d: douta_buf <= 22'h0000000000000000000000;
                12'h0b7e: douta_buf <= 22'h0000000000000000000000;
                12'h0b7f: douta_buf <= 22'h0000000000000000000000;
                12'h0b80: douta_buf <= 22'h0000000000000000000000;
                12'h0b81: douta_buf <= 22'h0000000000000000000000;
                12'h0b82: douta_buf <= 22'h0000000000000000000000;
                12'h0b83: douta_buf <= 22'h0000000000000000000000;
                12'h0b84: douta_buf <= 22'h0000000000000000000000;
                12'h0b85: douta_buf <= 22'h0000000000000000000000;
                12'h0b86: douta_buf <= 22'h0000000000000000000000;
                12'h0b87: douta_buf <= 22'h0000000000000000000000;
                12'h0b88: douta_buf <= 22'h0000000000000000000000;
                12'h0b89: douta_buf <= 22'h0000000000000000000000;
                12'h0b8a: douta_buf <= 22'h0000000000000000000000;
                12'h0b8b: douta_buf <= 22'h0000000000000000000000;
                12'h0b8c: douta_buf <= 22'h0000000000000000000000;
                12'h0b8d: douta_buf <= 22'h0000000000000000000000;
                12'h0b8e: douta_buf <= 22'h0000000000000000000000;
                12'h0b8f: douta_buf <= 22'h0000000000000000000000;
                12'h0b90: douta_buf <= 22'h0000000000000000000000;
                12'h0b91: douta_buf <= 22'h0000000000000000000000;
                12'h0b92: douta_buf <= 22'h0000000000000000000000;
                12'h0b93: douta_buf <= 22'h0000000000000000000000;
                12'h0b94: douta_buf <= 22'h0000000000000000000000;
                12'h0b95: douta_buf <= 22'h0000000000000000000000;
                12'h0b96: douta_buf <= 22'h0000000000000000000000;
                12'h0b97: douta_buf <= 22'h0000000000000000000000;
                12'h0b98: douta_buf <= 22'h0000000000000000000000;
                12'h0b99: douta_buf <= 22'h0000000000000000000000;
                12'h0b9a: douta_buf <= 22'h0000000000000000000000;
                12'h0b9b: douta_buf <= 22'h0000000000000000000000;
                12'h0b9c: douta_buf <= 22'h0000000000000000000000;
                12'h0b9d: douta_buf <= 22'h0000000000000000000000;
                12'h0b9e: douta_buf <= 22'h0000000000000000000000;
                12'h0b9f: douta_buf <= 22'h0000000000000000000000;
                12'h0ba0: douta_buf <= 22'h0000000000000000000000;
                12'h0ba1: douta_buf <= 22'h0000000000000000000000;
                12'h0ba2: douta_buf <= 22'h0000000000000000000000;
                12'h0ba3: douta_buf <= 22'h0000000000000000000000;
                12'h0ba4: douta_buf <= 22'h0000000000000000000000;
                12'h0ba5: douta_buf <= 22'h0000000000000000000000;
                12'h0ba6: douta_buf <= 22'h0000000000000000000000;
                12'h0ba7: douta_buf <= 22'h0000000000000000000000;
                12'h0ba8: douta_buf <= 22'h0000000000000000000000;
                12'h0ba9: douta_buf <= 22'h0000000000000000000000;
                12'h0baa: douta_buf <= 22'h0000000000000000000000;
                12'h0bab: douta_buf <= 22'h0000000000000000000000;
                12'h0bac: douta_buf <= 22'h0000000000000000000000;
                12'h0bad: douta_buf <= 22'h0000000000000000000000;
                12'h0bae: douta_buf <= 22'h0000000000000000000000;
                12'h0baf: douta_buf <= 22'h0000000000000000000000;
                12'h0bb0: douta_buf <= 22'h0000000000000000000000;
                12'h0bb1: douta_buf <= 22'h0000000000000000000000;
                12'h0bb2: douta_buf <= 22'h0000000000000000000000;
                12'h0bb3: douta_buf <= 22'h0000000000000000000000;
                12'h0bb4: douta_buf <= 22'h0000000000000000000000;
                12'h0bb5: douta_buf <= 22'h0000000000000000000000;
                12'h0bb6: douta_buf <= 22'h0000000000000000000000;
                12'h0bb7: douta_buf <= 22'h0000000000000000000000;
                12'h0bb8: douta_buf <= 22'h0000000000000000000000;
                12'h0bb9: douta_buf <= 22'h0000000000000000000000;
                12'h0bba: douta_buf <= 22'h0000000000000000000000;
                12'h0bbb: douta_buf <= 22'h0000000000000000000000;
                12'h0bbc: douta_buf <= 22'h0000000000000000000000;
                12'h0bbd: douta_buf <= 22'h0000000000000000000000;
                12'h0bbe: douta_buf <= 22'h0000000000000000000000;
                12'h0bbf: douta_buf <= 22'h0000000000000000000000;
                12'h0bc0: douta_buf <= 22'h0000000000000000000000;
                12'h0bc1: douta_buf <= 22'h0000000000000000000000;
                12'h0bc2: douta_buf <= 22'h0000000000000000000000;
                12'h0bc3: douta_buf <= 22'h0000000000000000000000;
                12'h0bc4: douta_buf <= 22'h0000000000000000000000;
                12'h0bc5: douta_buf <= 22'h0000000000000000000000;
                12'h0bc6: douta_buf <= 22'h0000000000000000000000;
                12'h0bc7: douta_buf <= 22'h0000000000000000000000;
                12'h0bc8: douta_buf <= 22'h0000000000000000000000;
                12'h0bc9: douta_buf <= 22'h0000000000000000000000;
                12'h0bca: douta_buf <= 22'h0000000000000000000000;
                12'h0bcb: douta_buf <= 22'h0000000000000000000000;
                12'h0bcc: douta_buf <= 22'h0000000000000000000000;
                12'h0bcd: douta_buf <= 22'h0000000000000000000000;
                12'h0bce: douta_buf <= 22'h0000000000000000000000;
                12'h0bcf: douta_buf <= 22'h0000000000000000000000;
                12'h0bd0: douta_buf <= 22'h0000000000000000000000;
                12'h0bd1: douta_buf <= 22'h0000000000000000000000;
                12'h0bd2: douta_buf <= 22'h0000000000000000000000;
                12'h0bd3: douta_buf <= 22'h0000000000000000000000;
                12'h0bd4: douta_buf <= 22'h0000000000000000000000;
                12'h0bd5: douta_buf <= 22'h0000000000000000000000;
                12'h0bd6: douta_buf <= 22'h0000000000000000000000;
                12'h0bd7: douta_buf <= 22'h0000000000000000000000;
                12'h0bd8: douta_buf <= 22'h0000000000000000000000;
                12'h0bd9: douta_buf <= 22'h0000000000000000000000;
                12'h0bda: douta_buf <= 22'h0000000000000000000000;
                12'h0bdb: douta_buf <= 22'h0000000000000000000000;
                12'h0bdc: douta_buf <= 22'h0000000000000000000000;
                12'h0bdd: douta_buf <= 22'h0000000000000000000000;
                12'h0bde: douta_buf <= 22'h0000000000000000000000;
                12'h0bdf: douta_buf <= 22'h0000000000000000000000;
                12'h0be0: douta_buf <= 22'h0000000000000000000000;
                12'h0be1: douta_buf <= 22'h0000000000000000000000;
                12'h0be2: douta_buf <= 22'h0000000000000000000000;
                12'h0be3: douta_buf <= 22'h0000000000000000000000;
                12'h0be4: douta_buf <= 22'h0000000000000000000000;
                12'h0be5: douta_buf <= 22'h0000000000000000000000;
                12'h0be6: douta_buf <= 22'h0000000000000000000000;
                12'h0be7: douta_buf <= 22'h0000000000000000000000;
                12'h0be8: douta_buf <= 22'h0000000000000000000000;
                12'h0be9: douta_buf <= 22'h0000000000000000000000;
                12'h0bea: douta_buf <= 22'h0000000000000000000000;
                12'h0beb: douta_buf <= 22'h0000000000000000000000;
                12'h0bec: douta_buf <= 22'h0000000000000000000000;
                12'h0bed: douta_buf <= 22'h0000000000000000000000;
                12'h0bee: douta_buf <= 22'h0000000000000000000000;
                12'h0bef: douta_buf <= 22'h0000000000000000000000;
                12'h0bf0: douta_buf <= 22'h0000000000000000000000;
                12'h0bf1: douta_buf <= 22'h0000000000000000000000;
                12'h0bf2: douta_buf <= 22'h0000000000000000000000;
                12'h0bf3: douta_buf <= 22'h0000000000000000000000;
                12'h0bf4: douta_buf <= 22'h0000000000000000000000;
                12'h0bf5: douta_buf <= 22'h0000000000000000000000;
                12'h0bf6: douta_buf <= 22'h0000000000000000000000;
                12'h0bf7: douta_buf <= 22'h0000000000000000000000;
                12'h0bf8: douta_buf <= 22'h0000000000000000000000;
                12'h0bf9: douta_buf <= 22'h0000000000000000000000;
                12'h0bfa: douta_buf <= 22'h0000000000000000000000;
                12'h0bfb: douta_buf <= 22'h0000000000000000000000;
                12'h0bfc: douta_buf <= 22'h0000000000000000000000;
                12'h0bfd: douta_buf <= 22'h0000000000000000000000;
                12'h0bfe: douta_buf <= 22'h0000000000000000000000;
                12'h0bff: douta_buf <= 22'h0000000000000000000000;
                12'h0c00: douta_buf <= 22'h0000000000000000000000;
                12'h0c01: douta_buf <= 22'h0000000000000000000000;
                12'h0c02: douta_buf <= 22'h0000000000000000000000;
                12'h0c03: douta_buf <= 22'h0000000000000000000000;
                12'h0c04: douta_buf <= 22'h0000000000000000000000;
                12'h0c05: douta_buf <= 22'h0000000000000000000000;
                12'h0c06: douta_buf <= 22'h0000000000000000000000;
                12'h0c07: douta_buf <= 22'h0000000000000000000000;
                12'h0c08: douta_buf <= 22'h0000000000000000000000;
                12'h0c09: douta_buf <= 22'h0000000000000000000000;
                12'h0c0a: douta_buf <= 22'h0000000000000000000000;
                12'h0c0b: douta_buf <= 22'h0000000000000000000000;
                12'h0c0c: douta_buf <= 22'h0000000000000000000000;
                12'h0c0d: douta_buf <= 22'h0000000000000000000000;
                12'h0c0e: douta_buf <= 22'h0000000000000000000000;
                12'h0c0f: douta_buf <= 22'h0000000000000000000000;
                12'h0c10: douta_buf <= 22'h0000000000000000000000;
                12'h0c11: douta_buf <= 22'h0000000000000000000000;
                12'h0c12: douta_buf <= 22'h0000000000000000000000;
                12'h0c13: douta_buf <= 22'h0000000000000000000000;
                12'h0c14: douta_buf <= 22'h0000000000000000000000;
                12'h0c15: douta_buf <= 22'h0000000000000000000000;
                12'h0c16: douta_buf <= 22'h0000000000000000000000;
                12'h0c17: douta_buf <= 22'h0000000000000000000000;
                12'h0c18: douta_buf <= 22'h0000000000000000000000;
                12'h0c19: douta_buf <= 22'h0000000000000000000000;
                12'h0c1a: douta_buf <= 22'h0000000000000000000000;
                12'h0c1b: douta_buf <= 22'h0000000000000000000000;
                12'h0c1c: douta_buf <= 22'h0000000000000000000000;
                12'h0c1d: douta_buf <= 22'h0000000000000000000000;
                12'h0c1e: douta_buf <= 22'h0000000000000000000000;
                12'h0c1f: douta_buf <= 22'h0000000000000000000000;
                12'h0c20: douta_buf <= 22'h0000000000000000000000;
                12'h0c21: douta_buf <= 22'h0000000000000000000000;
                12'h0c22: douta_buf <= 22'h0000000000000000000000;
                12'h0c23: douta_buf <= 22'h0000000000000000000000;
                12'h0c24: douta_buf <= 22'h0000000000000000000000;
                12'h0c25: douta_buf <= 22'h0000000000000000000000;
                12'h0c26: douta_buf <= 22'h0000000000000000000000;
                12'h0c27: douta_buf <= 22'h0000000000000000000000;
                12'h0c28: douta_buf <= 22'h0000000000000000000000;
                12'h0c29: douta_buf <= 22'h0000000000000000000000;
                12'h0c2a: douta_buf <= 22'h0000000000000000000000;
                12'h0c2b: douta_buf <= 22'h0000000000000000000000;
                12'h0c2c: douta_buf <= 22'h0000000000000000000000;
                12'h0c2d: douta_buf <= 22'h0000000000000000000000;
                12'h0c2e: douta_buf <= 22'h0000000000000000000000;
                12'h0c2f: douta_buf <= 22'h0000000000000000000000;
                12'h0c30: douta_buf <= 22'h0000000000000000000000;
                12'h0c31: douta_buf <= 22'h0000000000000000000000;
                12'h0c32: douta_buf <= 22'h0000000000000000000000;
                12'h0c33: douta_buf <= 22'h0000000000000000000000;
                12'h0c34: douta_buf <= 22'h0000000000000000000000;
                12'h0c35: douta_buf <= 22'h0000000000000000000000;
                12'h0c36: douta_buf <= 22'h0000000000000000000000;
                12'h0c37: douta_buf <= 22'h0000000000000000000000;
                12'h0c38: douta_buf <= 22'h0000000000000000000000;
                12'h0c39: douta_buf <= 22'h0000000000000000000000;
                12'h0c3a: douta_buf <= 22'h0000000000000000000000;
                12'h0c3b: douta_buf <= 22'h0000000000000000000000;
                12'h0c3c: douta_buf <= 22'h0000000000000000000000;
                12'h0c3d: douta_buf <= 22'h0000000000000000000000;
                12'h0c3e: douta_buf <= 22'h0000000000000000000000;
                12'h0c3f: douta_buf <= 22'h0000000000000000000000;
                12'h0c40: douta_buf <= 22'h0000000000000000000000;
                12'h0c41: douta_buf <= 22'h0000000000000000000000;
                12'h0c42: douta_buf <= 22'h0000000000000000000000;
                12'h0c43: douta_buf <= 22'h0000000000000000000000;
                12'h0c44: douta_buf <= 22'h0000000000000000000000;
                12'h0c45: douta_buf <= 22'h0000000000000000000000;
                12'h0c46: douta_buf <= 22'h0000000000000000000000;
                12'h0c47: douta_buf <= 22'h0000000000000000000000;
                12'h0c48: douta_buf <= 22'h0000000000000000000000;
                12'h0c49: douta_buf <= 22'h0000000000000000000000;
                12'h0c4a: douta_buf <= 22'h0000000000000000000000;
                12'h0c4b: douta_buf <= 22'h0000000000000000000000;
                12'h0c4c: douta_buf <= 22'h0000000000000000000000;
                12'h0c4d: douta_buf <= 22'h0000000000000000000000;
                12'h0c4e: douta_buf <= 22'h0000000000000000000000;
                12'h0c4f: douta_buf <= 22'h0000000000000000000000;
                12'h0c50: douta_buf <= 22'h0000000000000000000000;
                12'h0c51: douta_buf <= 22'h0000000000000000000000;
                12'h0c52: douta_buf <= 22'h0000000000000000000000;
                12'h0c53: douta_buf <= 22'h0000000000000000000000;
                12'h0c54: douta_buf <= 22'h0000000000000000000000;
                12'h0c55: douta_buf <= 22'h0000000000000000000000;
                12'h0c56: douta_buf <= 22'h0000000000000000000000;
                12'h0c57: douta_buf <= 22'h0000000000000000000000;
                12'h0c58: douta_buf <= 22'h0000000000000000000000;
                12'h0c59: douta_buf <= 22'h0000000000000000000000;
                12'h0c5a: douta_buf <= 22'h0000000000000000000000;
                12'h0c5b: douta_buf <= 22'h0000000000000000000000;
                12'h0c5c: douta_buf <= 22'h0000000000000000000000;
                12'h0c5d: douta_buf <= 22'h0000000000000000000000;
                12'h0c5e: douta_buf <= 22'h0000000000000000000000;
                12'h0c5f: douta_buf <= 22'h0000000000000000000000;
                12'h0c60: douta_buf <= 22'h0000000000000000000000;
                12'h0c61: douta_buf <= 22'h0000000000000000000000;
                12'h0c62: douta_buf <= 22'h0000000000000000000000;
                12'h0c63: douta_buf <= 22'h0000000000000000000000;
                12'h0c64: douta_buf <= 22'h0000000000000000000000;
                12'h0c65: douta_buf <= 22'h0000000000000000000000;
                12'h0c66: douta_buf <= 22'h0000000000000000000000;
                12'h0c67: douta_buf <= 22'h0000000000000000000000;
                12'h0c68: douta_buf <= 22'h0000000000000000000000;
                12'h0c69: douta_buf <= 22'h0000000000000000000000;
                12'h0c6a: douta_buf <= 22'h0000000000000000000000;
                12'h0c6b: douta_buf <= 22'h0000000000000000000000;
                12'h0c6c: douta_buf <= 22'h0000000000000000000000;
                12'h0c6d: douta_buf <= 22'h0000000000000000000000;
                12'h0c6e: douta_buf <= 22'h0000000000000000000000;
                12'h0c6f: douta_buf <= 22'h0000000000000000000000;
                12'h0c70: douta_buf <= 22'h0000000000000000000000;
                12'h0c71: douta_buf <= 22'h0000000000000000000000;
                12'h0c72: douta_buf <= 22'h0000000000000000000000;
                12'h0c73: douta_buf <= 22'h0000000000000000000000;
                12'h0c74: douta_buf <= 22'h0000000000000000000000;
                12'h0c75: douta_buf <= 22'h0000000000000000000000;
                12'h0c76: douta_buf <= 22'h0000000000000000000000;
                12'h0c77: douta_buf <= 22'h0000000000000000000000;
                12'h0c78: douta_buf <= 22'h0000000000000000000000;
                12'h0c79: douta_buf <= 22'h0000000000000000000000;
                12'h0c7a: douta_buf <= 22'h0000000000000000000000;
                12'h0c7b: douta_buf <= 22'h0000000000000000000000;
                12'h0c7c: douta_buf <= 22'h0000000000000000000000;
                12'h0c7d: douta_buf <= 22'h0000000000000000000000;
                12'h0c7e: douta_buf <= 22'h0000000000000000000000;
                12'h0c7f: douta_buf <= 22'h0000000000000000000000;
                12'h0c80: douta_buf <= 22'h0000000000000000000000;
                12'h0c81: douta_buf <= 22'h0000000000000000000000;
                12'h0c82: douta_buf <= 22'h0000000000000000000000;
                12'h0c83: douta_buf <= 22'h0000000000000000000000;
                12'h0c84: douta_buf <= 22'h0000000000000000000000;
                12'h0c85: douta_buf <= 22'h0000000000000000000000;
                12'h0c86: douta_buf <= 22'h0000000000000000000000;
                12'h0c87: douta_buf <= 22'h0000000000000000000000;
                12'h0c88: douta_buf <= 22'h0000000000000000000000;
                12'h0c89: douta_buf <= 22'h0000000000000000000000;
                12'h0c8a: douta_buf <= 22'h0000000000000000000000;
                12'h0c8b: douta_buf <= 22'h0000000000000000000000;
                12'h0c8c: douta_buf <= 22'h0000000000000000000000;
                12'h0c8d: douta_buf <= 22'h0000000000000000000000;
                12'h0c8e: douta_buf <= 22'h0000000000000000000000;
                12'h0c8f: douta_buf <= 22'h0000000000000000000000;
                12'h0c90: douta_buf <= 22'h0000000000000000000000;
                12'h0c91: douta_buf <= 22'h0000000000000000000000;
                12'h0c92: douta_buf <= 22'h0000000000000000000000;
                12'h0c93: douta_buf <= 22'h0000000000000000000000;
                12'h0c94: douta_buf <= 22'h0000000000000000000000;
                12'h0c95: douta_buf <= 22'h0000000000000000000000;
                12'h0c96: douta_buf <= 22'h0000000000000000000000;
                12'h0c97: douta_buf <= 22'h0000000000000000000000;
                12'h0c98: douta_buf <= 22'h0000000000000000000000;
                12'h0c99: douta_buf <= 22'h0000000000000000000000;
                12'h0c9a: douta_buf <= 22'h0000000000000000000000;
                12'h0c9b: douta_buf <= 22'h0000000000000000000000;
                12'h0c9c: douta_buf <= 22'h0000000000000000000000;
                12'h0c9d: douta_buf <= 22'h0000000000000000000000;
                12'h0c9e: douta_buf <= 22'h0000000000000000000000;
                12'h0c9f: douta_buf <= 22'h0000000000000000000000;
                12'h0ca0: douta_buf <= 22'h0000000000000000000000;
                12'h0ca1: douta_buf <= 22'h0000000000000000000000;
                12'h0ca2: douta_buf <= 22'h0000000000000000000000;
                12'h0ca3: douta_buf <= 22'h0000000000000000000000;
                12'h0ca4: douta_buf <= 22'h0000000000000000000000;
                12'h0ca5: douta_buf <= 22'h0000000000000000000000;
                12'h0ca6: douta_buf <= 22'h0000000000000000000000;
                12'h0ca7: douta_buf <= 22'h0000000000000000000000;
                12'h0ca8: douta_buf <= 22'h0000000000000000000000;
                12'h0ca9: douta_buf <= 22'h0000000000000000000000;
                12'h0caa: douta_buf <= 22'h0000000000000000000000;
                12'h0cab: douta_buf <= 22'h0000000000000000000000;
                12'h0cac: douta_buf <= 22'h0000000000000000000000;
                12'h0cad: douta_buf <= 22'h0000000000000000000000;
                12'h0cae: douta_buf <= 22'h0000000000000000000000;
                12'h0caf: douta_buf <= 22'h0000000000000000000000;
                12'h0cb0: douta_buf <= 22'h0000000000000000000000;
                12'h0cb1: douta_buf <= 22'h0000000000000000000000;
                12'h0cb2: douta_buf <= 22'h0000000000000000000000;
                12'h0cb3: douta_buf <= 22'h0000000000000000000000;
                12'h0cb4: douta_buf <= 22'h0000000000000000000000;
                12'h0cb5: douta_buf <= 22'h0000000000000000000000;
                12'h0cb6: douta_buf <= 22'h0000000000000000000000;
                12'h0cb7: douta_buf <= 22'h0000000000000000000000;
                12'h0cb8: douta_buf <= 22'h0000000000000000000000;
                12'h0cb9: douta_buf <= 22'h0000000000000000000000;
                12'h0cba: douta_buf <= 22'h0000000000000000000000;
                12'h0cbb: douta_buf <= 22'h0000000000000000000000;
                12'h0cbc: douta_buf <= 22'h0000000000000000000000;
                12'h0cbd: douta_buf <= 22'h0000000000000000000000;
                12'h0cbe: douta_buf <= 22'h0000000000000000000000;
                12'h0cbf: douta_buf <= 22'h0000000000000000000000;
                12'h0cc0: douta_buf <= 22'h0000000000000000000000;
                12'h0cc1: douta_buf <= 22'h0000000000000000000000;
                12'h0cc2: douta_buf <= 22'h0000000000000000000000;
                12'h0cc3: douta_buf <= 22'h0000000000000000000000;
                12'h0cc4: douta_buf <= 22'h0000000000000000000000;
                12'h0cc5: douta_buf <= 22'h0000000000000000000000;
                12'h0cc6: douta_buf <= 22'h0000000000000000000000;
                12'h0cc7: douta_buf <= 22'h0000000000000000000000;
                12'h0cc8: douta_buf <= 22'h0000000000000000000000;
                12'h0cc9: douta_buf <= 22'h0000000000000000000000;
                12'h0cca: douta_buf <= 22'h0000000000000000000000;
                12'h0ccb: douta_buf <= 22'h0000000000000000000000;
                12'h0ccc: douta_buf <= 22'h0000000000000000000000;
                12'h0ccd: douta_buf <= 22'h0000000000000000000000;
                12'h0cce: douta_buf <= 22'h0000000000000000000000;
                12'h0ccf: douta_buf <= 22'h0000000000000000000000;
                12'h0cd0: douta_buf <= 22'h0000000000000000000000;
                12'h0cd1: douta_buf <= 22'h0000000000000000000000;
                12'h0cd2: douta_buf <= 22'h0000000000000000000000;
                12'h0cd3: douta_buf <= 22'h0000000000000000000000;
                12'h0cd4: douta_buf <= 22'h0000000000000000000000;
                12'h0cd5: douta_buf <= 22'h0000000000000000000000;
                12'h0cd6: douta_buf <= 22'h0000000000000000000000;
                12'h0cd7: douta_buf <= 22'h0000000000000000000000;
                12'h0cd8: douta_buf <= 22'h0000000000000000000000;
                12'h0cd9: douta_buf <= 22'h0000000000000000000000;
                12'h0cda: douta_buf <= 22'h0000000000000000000000;
                12'h0cdb: douta_buf <= 22'h0000000000000000000000;
                12'h0cdc: douta_buf <= 22'h0000000000000000000000;
                12'h0cdd: douta_buf <= 22'h0000000000000000000000;
                12'h0cde: douta_buf <= 22'h0000000000000000000000;
                12'h0cdf: douta_buf <= 22'h0000000000000000000000;
                12'h0ce0: douta_buf <= 22'h0000000000000000000000;
                12'h0ce1: douta_buf <= 22'h0000000000000000000000;
                12'h0ce2: douta_buf <= 22'h0000000000000000000000;
                12'h0ce3: douta_buf <= 22'h0000000000000000000000;
                12'h0ce4: douta_buf <= 22'h0000000000000000000000;
                12'h0ce5: douta_buf <= 22'h0000000000000000000000;
                12'h0ce6: douta_buf <= 22'h0000000000000000000000;
                12'h0ce7: douta_buf <= 22'h0000000000000000000000;
                12'h0ce8: douta_buf <= 22'h0000000000000000000000;
                12'h0ce9: douta_buf <= 22'h0000000000000000000000;
                12'h0cea: douta_buf <= 22'h0000000000000000000000;
                12'h0ceb: douta_buf <= 22'h0000000000000000000000;
                12'h0cec: douta_buf <= 22'h0000000000000000000000;
                12'h0ced: douta_buf <= 22'h0000000000000000000000;
                12'h0cee: douta_buf <= 22'h0000000000000000000000;
                12'h0cef: douta_buf <= 22'h0000000000000000000000;
                12'h0cf0: douta_buf <= 22'h0000000000000000000000;
                12'h0cf1: douta_buf <= 22'h0000000000000000000000;
                12'h0cf2: douta_buf <= 22'h0000000000000000000000;
                12'h0cf3: douta_buf <= 22'h0000000000000000000000;
                12'h0cf4: douta_buf <= 22'h0000000000000000000000;
                12'h0cf5: douta_buf <= 22'h0000000000000000000000;
                12'h0cf6: douta_buf <= 22'h0000000000000000000000;
                12'h0cf7: douta_buf <= 22'h0000000000000000000000;
                12'h0cf8: douta_buf <= 22'h0000000000000000000000;
                12'h0cf9: douta_buf <= 22'h0000000000000000000000;
                12'h0cfa: douta_buf <= 22'h0000000000000000000000;
                12'h0cfb: douta_buf <= 22'h0000000000000000000000;
                12'h0cfc: douta_buf <= 22'h0000000000000000000000;
                12'h0cfd: douta_buf <= 22'h0000000000000000000000;
                12'h0cfe: douta_buf <= 22'h0000000000000000000000;
                12'h0cff: douta_buf <= 22'h0000000000000000000000;
                12'h0d00: douta_buf <= 22'h0000000000000000000000;
                12'h0d01: douta_buf <= 22'h0000000000000000000000;
                12'h0d02: douta_buf <= 22'h0000000000000000000000;
                12'h0d03: douta_buf <= 22'h0000000000000000000000;
                12'h0d04: douta_buf <= 22'h0000000000000000000000;
                12'h0d05: douta_buf <= 22'h0000000000000000000000;
                12'h0d06: douta_buf <= 22'h0000000000000000000000;
                12'h0d07: douta_buf <= 22'h0000000000000000000000;
                12'h0d08: douta_buf <= 22'h0000000000000000000000;
                12'h0d09: douta_buf <= 22'h0000000000000000000000;
                12'h0d0a: douta_buf <= 22'h0000000000000000000000;
                12'h0d0b: douta_buf <= 22'h0000000000000000000000;
                12'h0d0c: douta_buf <= 22'h0000000000000000000000;
                12'h0d0d: douta_buf <= 22'h0000000000000000000000;
                12'h0d0e: douta_buf <= 22'h0000000000000000000000;
                12'h0d0f: douta_buf <= 22'h0000000000000000000000;
                12'h0d10: douta_buf <= 22'h0000000000000000000000;
                12'h0d11: douta_buf <= 22'h0000000000000000000000;
                12'h0d12: douta_buf <= 22'h0000000000000000000000;
                12'h0d13: douta_buf <= 22'h0000000000000000000000;
                12'h0d14: douta_buf <= 22'h0000000000000000000000;
                12'h0d15: douta_buf <= 22'h0000000000000000000000;
                12'h0d16: douta_buf <= 22'h0000000000000000000000;
                12'h0d17: douta_buf <= 22'h0000000000000000000000;
                12'h0d18: douta_buf <= 22'h0000000000000000000000;
                12'h0d19: douta_buf <= 22'h0000000000000000000000;
                12'h0d1a: douta_buf <= 22'h0000000000000000000000;
                12'h0d1b: douta_buf <= 22'h0000000000000000000000;
                12'h0d1c: douta_buf <= 22'h0000000000000000000000;
                12'h0d1d: douta_buf <= 22'h0000000000000000000000;
                12'h0d1e: douta_buf <= 22'h0000000000000000000000;
                12'h0d1f: douta_buf <= 22'h0000000000000000000000;
                12'h0d20: douta_buf <= 22'h0000000000000000000000;
                12'h0d21: douta_buf <= 22'h0000000000000000000000;
                12'h0d22: douta_buf <= 22'h0000000000000000000000;
                12'h0d23: douta_buf <= 22'h0000000000000000000000;
                12'h0d24: douta_buf <= 22'h0000000000000000000000;
                12'h0d25: douta_buf <= 22'h0000000000000000000000;
                12'h0d26: douta_buf <= 22'h0000000000000000000000;
                12'h0d27: douta_buf <= 22'h0000000000000000000000;
                12'h0d28: douta_buf <= 22'h0000000000000000000000;
                12'h0d29: douta_buf <= 22'h0000000000000000000000;
                12'h0d2a: douta_buf <= 22'h0000000000000000000000;
                12'h0d2b: douta_buf <= 22'h0000000000000000000000;
                12'h0d2c: douta_buf <= 22'h0000000000000000000000;
                12'h0d2d: douta_buf <= 22'h0000000000000000000000;
                12'h0d2e: douta_buf <= 22'h0000000000000000000000;
                12'h0d2f: douta_buf <= 22'h0000000000000000000000;
                12'h0d30: douta_buf <= 22'h0000000000000000000000;
                12'h0d31: douta_buf <= 22'h0000000000000000000000;
                12'h0d32: douta_buf <= 22'h0000000000000000000000;
                12'h0d33: douta_buf <= 22'h0000000000000000000000;
                12'h0d34: douta_buf <= 22'h0000000000000000000000;
                12'h0d35: douta_buf <= 22'h0000000000000000000000;
                12'h0d36: douta_buf <= 22'h0000000000000000000000;
                12'h0d37: douta_buf <= 22'h0000000000000000000000;
                12'h0d38: douta_buf <= 22'h0000000000000000000000;
                12'h0d39: douta_buf <= 22'h0000000000000000000000;
                12'h0d3a: douta_buf <= 22'h0000000000000000000000;
                12'h0d3b: douta_buf <= 22'h0000000000000000000000;
                12'h0d3c: douta_buf <= 22'h0000000000000000000000;
                12'h0d3d: douta_buf <= 22'h0000000000000000000000;
                12'h0d3e: douta_buf <= 22'h0000000000000000000000;
                12'h0d3f: douta_buf <= 22'h0000000000000000000000;
                12'h0d40: douta_buf <= 22'h0000000000000000000000;
                12'h0d41: douta_buf <= 22'h0000000000000000000000;
                12'h0d42: douta_buf <= 22'h0000000000000000000000;
                12'h0d43: douta_buf <= 22'h0000000000000000000000;
                12'h0d44: douta_buf <= 22'h0000000000000000000000;
                12'h0d45: douta_buf <= 22'h0000000000000000000000;
                12'h0d46: douta_buf <= 22'h0000000000000000000000;
                12'h0d47: douta_buf <= 22'h0000000000000000000000;
                12'h0d48: douta_buf <= 22'h0000000000000000000000;
                12'h0d49: douta_buf <= 22'h0000000000000000000000;
                12'h0d4a: douta_buf <= 22'h0000000000000000000000;
                12'h0d4b: douta_buf <= 22'h0000000000000000000000;
                12'h0d4c: douta_buf <= 22'h0000000000000000000000;
                12'h0d4d: douta_buf <= 22'h0000000000000000000000;
                12'h0d4e: douta_buf <= 22'h0000000000000000000000;
                12'h0d4f: douta_buf <= 22'h0000000000000000000000;
                12'h0d50: douta_buf <= 22'h0000000000000000000000;
                12'h0d51: douta_buf <= 22'h0000000000000000000000;
                12'h0d52: douta_buf <= 22'h0000000000000000000000;
                12'h0d53: douta_buf <= 22'h0000000000000000000000;
                12'h0d54: douta_buf <= 22'h0000000000000000000000;
                12'h0d55: douta_buf <= 22'h0000000000000000000000;
                12'h0d56: douta_buf <= 22'h0000000000000000000000;
                12'h0d57: douta_buf <= 22'h0000000000000000000000;
                12'h0d58: douta_buf <= 22'h0000000000000000000000;
                12'h0d59: douta_buf <= 22'h0000000000000000000000;
                12'h0d5a: douta_buf <= 22'h0000000000000000000000;
                12'h0d5b: douta_buf <= 22'h0000000000000000000000;
                12'h0d5c: douta_buf <= 22'h0000000000000000000000;
                12'h0d5d: douta_buf <= 22'h0000000000000000000000;
                12'h0d5e: douta_buf <= 22'h0000000000000000000000;
                12'h0d5f: douta_buf <= 22'h0000000000000000000000;
                12'h0d60: douta_buf <= 22'h0000000000000000000000;
                12'h0d61: douta_buf <= 22'h0000000000000000000000;
                12'h0d62: douta_buf <= 22'h0000000000000000000000;
                12'h0d63: douta_buf <= 22'h0000000000000000000000;
                12'h0d64: douta_buf <= 22'h0000000000000000000000;
                12'h0d65: douta_buf <= 22'h0000000000000000000000;
                12'h0d66: douta_buf <= 22'h0000000000000000000000;
                12'h0d67: douta_buf <= 22'h0000000000000000000000;
                12'h0d68: douta_buf <= 22'h0000000000000000000000;
                12'h0d69: douta_buf <= 22'h0000000000000000000000;
                12'h0d6a: douta_buf <= 22'h0000000000000000000000;
                12'h0d6b: douta_buf <= 22'h0000000000000000000000;
                12'h0d6c: douta_buf <= 22'h0000000000000000000000;
                12'h0d6d: douta_buf <= 22'h0000000000000000000000;
                12'h0d6e: douta_buf <= 22'h0000000000000000000000;
                12'h0d6f: douta_buf <= 22'h0000000000000000000000;
                12'h0d70: douta_buf <= 22'h0000000000000000000000;
                12'h0d71: douta_buf <= 22'h0000000000000000000000;
                12'h0d72: douta_buf <= 22'h0000000000000000000000;
                12'h0d73: douta_buf <= 22'h0000000000000000000000;
                12'h0d74: douta_buf <= 22'h0000000000000000000000;
                12'h0d75: douta_buf <= 22'h0000000000000000000000;
                12'h0d76: douta_buf <= 22'h0000000000000000000000;
                12'h0d77: douta_buf <= 22'h0000000000000000000000;
                12'h0d78: douta_buf <= 22'h0000000000000000000000;
                12'h0d79: douta_buf <= 22'h0000000000000000000000;
                12'h0d7a: douta_buf <= 22'h0000000000000000000000;
                12'h0d7b: douta_buf <= 22'h0000000000000000000000;
                12'h0d7c: douta_buf <= 22'h0000000000000000000000;
                12'h0d7d: douta_buf <= 22'h0000000000000000000000;
                12'h0d7e: douta_buf <= 22'h0000000000000000000000;
                12'h0d7f: douta_buf <= 22'h0000000000000000000000;
                12'h0d80: douta_buf <= 22'h0000000000000000000000;
                12'h0d81: douta_buf <= 22'h0000000000000000000000;
                12'h0d82: douta_buf <= 22'h0000000000000000000000;
                12'h0d83: douta_buf <= 22'h0000000000000000000000;
                12'h0d84: douta_buf <= 22'h0000000000000000000000;
                12'h0d85: douta_buf <= 22'h0000000000000000000000;
                12'h0d86: douta_buf <= 22'h0000000000000000000000;
                12'h0d87: douta_buf <= 22'h0000000000000000000000;
                12'h0d88: douta_buf <= 22'h0000000000000000000000;
                12'h0d89: douta_buf <= 22'h0000000000000000000000;
                12'h0d8a: douta_buf <= 22'h0000000000000000000000;
                12'h0d8b: douta_buf <= 22'h0000000000000000000000;
                12'h0d8c: douta_buf <= 22'h0000000000000000000000;
                12'h0d8d: douta_buf <= 22'h0000000000000000000000;
                12'h0d8e: douta_buf <= 22'h0000000000000000000000;
                12'h0d8f: douta_buf <= 22'h0000000000000000000000;
                12'h0d90: douta_buf <= 22'h0000000000000000000000;
                12'h0d91: douta_buf <= 22'h0000000000000000000000;
                12'h0d92: douta_buf <= 22'h0000000000000000000000;
                12'h0d93: douta_buf <= 22'h0000000000000000000000;
                12'h0d94: douta_buf <= 22'h0000000000000000000000;
                12'h0d95: douta_buf <= 22'h0000000000000000000000;
                12'h0d96: douta_buf <= 22'h0000000000000000000000;
                12'h0d97: douta_buf <= 22'h0000000000000000000000;
                12'h0d98: douta_buf <= 22'h0000000000000000000000;
                12'h0d99: douta_buf <= 22'h0000000000000000000000;
                12'h0d9a: douta_buf <= 22'h0000000000000000000000;
                12'h0d9b: douta_buf <= 22'h0000000000000000000000;
                12'h0d9c: douta_buf <= 22'h0000000000000000000000;
                12'h0d9d: douta_buf <= 22'h0000000000000000000000;
                12'h0d9e: douta_buf <= 22'h0000000000000000000000;
                12'h0d9f: douta_buf <= 22'h0000000000000000000000;
                12'h0da0: douta_buf <= 22'h0000000000000000000000;
                12'h0da1: douta_buf <= 22'h0000000000000000000000;
                12'h0da2: douta_buf <= 22'h0000000000000000000000;
                12'h0da3: douta_buf <= 22'h0000000000000000000000;
                12'h0da4: douta_buf <= 22'h0000000000000000000000;
                12'h0da5: douta_buf <= 22'h0000000000000000000000;
                12'h0da6: douta_buf <= 22'h0000000000000000000000;
                12'h0da7: douta_buf <= 22'h0000000000000000000000;
                12'h0da8: douta_buf <= 22'h0000000000000000000000;
                12'h0da9: douta_buf <= 22'h0000000000000000000000;
                12'h0daa: douta_buf <= 22'h0000000000000000000000;
                12'h0dab: douta_buf <= 22'h0000000000000000000000;
                12'h0dac: douta_buf <= 22'h0000000000000000000000;
                12'h0dad: douta_buf <= 22'h0000000000000000000000;
                12'h0dae: douta_buf <= 22'h0000000000000000000000;
                12'h0daf: douta_buf <= 22'h0000000000000000000000;
                12'h0db0: douta_buf <= 22'h0000000000000000000000;
                12'h0db1: douta_buf <= 22'h0000000000000000000000;
                12'h0db2: douta_buf <= 22'h0000000000000000000000;
                12'h0db3: douta_buf <= 22'h0000000000000000000000;
                12'h0db4: douta_buf <= 22'h0000000000000000000000;
                12'h0db5: douta_buf <= 22'h0000000000000000000000;
                12'h0db6: douta_buf <= 22'h0000000000000000000000;
                12'h0db7: douta_buf <= 22'h0000000000000000000000;
                12'h0db8: douta_buf <= 22'h0000000000000000000000;
                12'h0db9: douta_buf <= 22'h0000000000000000000000;
                12'h0dba: douta_buf <= 22'h0000000000000000000000;
                12'h0dbb: douta_buf <= 22'h0000000000000000000000;
                12'h0dbc: douta_buf <= 22'h0000000000000000000000;
                12'h0dbd: douta_buf <= 22'h0000000000000000000000;
                12'h0dbe: douta_buf <= 22'h0000000000000000000000;
                12'h0dbf: douta_buf <= 22'h0000000000000000000000;
                12'h0dc0: douta_buf <= 22'h0000000000000000000000;
                12'h0dc1: douta_buf <= 22'h0000000000000000000000;
                12'h0dc2: douta_buf <= 22'h0000000000000000000000;
                12'h0dc3: douta_buf <= 22'h0000000000000000000000;
                12'h0dc4: douta_buf <= 22'h0000000000000000000000;
                12'h0dc5: douta_buf <= 22'h0000000000000000000000;
                12'h0dc6: douta_buf <= 22'h0000000000000000000000;
                12'h0dc7: douta_buf <= 22'h0000000000000000000000;
                12'h0dc8: douta_buf <= 22'h0000000000000000000000;
                12'h0dc9: douta_buf <= 22'h0000000000000000000000;
                12'h0dca: douta_buf <= 22'h0000000000000000000000;
                12'h0dcb: douta_buf <= 22'h0000000000000000000000;
                12'h0dcc: douta_buf <= 22'h0000000000000000000000;
                12'h0dcd: douta_buf <= 22'h0000000000000000000000;
                12'h0dce: douta_buf <= 22'h0000000000000000000000;
                12'h0dcf: douta_buf <= 22'h0000000000000000000000;
                12'h0dd0: douta_buf <= 22'h0000000000000000000000;
                12'h0dd1: douta_buf <= 22'h0000000000000000000000;
                12'h0dd2: douta_buf <= 22'h0000000000000000000000;
                12'h0dd3: douta_buf <= 22'h0000000000000000000000;
                12'h0dd4: douta_buf <= 22'h0000000000000000000000;
                12'h0dd5: douta_buf <= 22'h0000000000000000000000;
                12'h0dd6: douta_buf <= 22'h0000000000000000000000;
                12'h0dd7: douta_buf <= 22'h0000000000000000000000;
                12'h0dd8: douta_buf <= 22'h0000000000000000000000;
                12'h0dd9: douta_buf <= 22'h0000000000000000000000;
                12'h0dda: douta_buf <= 22'h0000000000000000000000;
                12'h0ddb: douta_buf <= 22'h0000000000000000000000;
                12'h0ddc: douta_buf <= 22'h0000000000000000000000;
                12'h0ddd: douta_buf <= 22'h0000000000000000000000;
                12'h0dde: douta_buf <= 22'h0000000000000000000000;
                12'h0ddf: douta_buf <= 22'h0000000000000000000000;
                12'h0de0: douta_buf <= 22'h0000000000000000000000;
                12'h0de1: douta_buf <= 22'h0000000000000000000000;
                12'h0de2: douta_buf <= 22'h0000000000000000000000;
                12'h0de3: douta_buf <= 22'h0000000000000000000000;
                12'h0de4: douta_buf <= 22'h0000000000000000000000;
                12'h0de5: douta_buf <= 22'h0000000000000000000000;
                12'h0de6: douta_buf <= 22'h0000000000000000000000;
                12'h0de7: douta_buf <= 22'h0000000000000000000000;
                12'h0de8: douta_buf <= 22'h0000000000000000000000;
                12'h0de9: douta_buf <= 22'h0000000000000000000000;
                12'h0dea: douta_buf <= 22'h0000000000000000000000;
                12'h0deb: douta_buf <= 22'h0000000000000000000000;
                12'h0dec: douta_buf <= 22'h0000000000000000000000;
                12'h0ded: douta_buf <= 22'h0000000000000000000000;
                12'h0dee: douta_buf <= 22'h0000000000000000000000;
                12'h0def: douta_buf <= 22'h0000000000000000000000;
                12'h0df0: douta_buf <= 22'h0000000000000000000000;
                12'h0df1: douta_buf <= 22'h0000000000000000000000;
                12'h0df2: douta_buf <= 22'h0000000000000000000000;
                12'h0df3: douta_buf <= 22'h0000000000000000000000;
                12'h0df4: douta_buf <= 22'h0000000000000000000000;
                12'h0df5: douta_buf <= 22'h0000000000000000000000;
                12'h0df6: douta_buf <= 22'h0000000000000000000000;
                12'h0df7: douta_buf <= 22'h0000000000000000000000;
                12'h0df8: douta_buf <= 22'h0000000000000000000000;
                12'h0df9: douta_buf <= 22'h0000000000000000000000;
                12'h0dfa: douta_buf <= 22'h0000000000000000000000;
                12'h0dfb: douta_buf <= 22'h0000000000000000000000;
                12'h0dfc: douta_buf <= 22'h0000000000000000000000;
                12'h0dfd: douta_buf <= 22'h0000000000000000000000;
                12'h0dfe: douta_buf <= 22'h0000000000000000000000;
                12'h0dff: douta_buf <= 22'h0000000000000000000000;
                12'h0e00: douta_buf <= 22'h0000000000000000000000;
                12'h0e01: douta_buf <= 22'h0000000000000000000000;
                12'h0e02: douta_buf <= 22'h0000000000000000000000;
                12'h0e03: douta_buf <= 22'h0000000000000000000000;
                12'h0e04: douta_buf <= 22'h0000000000000000000000;
                12'h0e05: douta_buf <= 22'h0000000000000000000000;
                12'h0e06: douta_buf <= 22'h0000000000000000000000;
                12'h0e07: douta_buf <= 22'h0000000000000000000000;
                12'h0e08: douta_buf <= 22'h0000000000000000000000;
                12'h0e09: douta_buf <= 22'h0000000000000000000000;
                12'h0e0a: douta_buf <= 22'h0000000000000000000000;
                12'h0e0b: douta_buf <= 22'h0000000000000000000000;
                12'h0e0c: douta_buf <= 22'h0000000000000000000000;
                12'h0e0d: douta_buf <= 22'h0000000000000000000000;
                12'h0e0e: douta_buf <= 22'h0000000000000000000000;
                12'h0e0f: douta_buf <= 22'h0000000000000000000000;
                12'h0e10: douta_buf <= 22'h0000000000000000000000;
                12'h0e11: douta_buf <= 22'h0000000000000000000000;
                12'h0e12: douta_buf <= 22'h0000000000000000000000;
                12'h0e13: douta_buf <= 22'h0000000000000000000000;
                12'h0e14: douta_buf <= 22'h0000000000000000000000;
                12'h0e15: douta_buf <= 22'h0000000000000000000000;
                12'h0e16: douta_buf <= 22'h0000000000000000000000;
                12'h0e17: douta_buf <= 22'h0000000000000000000000;
                12'h0e18: douta_buf <= 22'h0000000000000000000000;
                12'h0e19: douta_buf <= 22'h0000000000000000000000;
                12'h0e1a: douta_buf <= 22'h0000000000000000000000;
                12'h0e1b: douta_buf <= 22'h0000000000000000000000;
                12'h0e1c: douta_buf <= 22'h0000000000000000000000;
                12'h0e1d: douta_buf <= 22'h0000000000000000000000;
                12'h0e1e: douta_buf <= 22'h0000000000000000000000;
                12'h0e1f: douta_buf <= 22'h0000000000000000000000;
                12'h0e20: douta_buf <= 22'h0000000000000000000000;
                12'h0e21: douta_buf <= 22'h0000000000000000000000;
                12'h0e22: douta_buf <= 22'h0000000000000000000000;
                12'h0e23: douta_buf <= 22'h0000000000000000000000;
                12'h0e24: douta_buf <= 22'h0000000000000000000000;
                12'h0e25: douta_buf <= 22'h0000000000000000000000;
                12'h0e26: douta_buf <= 22'h0000000000000000000000;
                12'h0e27: douta_buf <= 22'h0000000000000000000000;
                12'h0e28: douta_buf <= 22'h0000000000000000000000;
                12'h0e29: douta_buf <= 22'h0000000000000000000000;
                12'h0e2a: douta_buf <= 22'h0000000000000000000000;
                12'h0e2b: douta_buf <= 22'h0000000000000000000000;
                12'h0e2c: douta_buf <= 22'h0000000000000000000000;
                12'h0e2d: douta_buf <= 22'h0000000000000000000000;
                12'h0e2e: douta_buf <= 22'h0000000000000000000000;
                12'h0e2f: douta_buf <= 22'h0000000000000000000000;
                12'h0e30: douta_buf <= 22'h0000000000000000000000;
                12'h0e31: douta_buf <= 22'h0000000000000000000000;
                12'h0e32: douta_buf <= 22'h0000000000000000000000;
                12'h0e33: douta_buf <= 22'h0000000000000000000000;
                12'h0e34: douta_buf <= 22'h0000000000000000000000;
                12'h0e35: douta_buf <= 22'h0000000000000000000000;
                12'h0e36: douta_buf <= 22'h0000000000000000000000;
                12'h0e37: douta_buf <= 22'h0000000000000000000000;
                12'h0e38: douta_buf <= 22'h0000000000000000000000;
                12'h0e39: douta_buf <= 22'h0000000000000000000000;
                12'h0e3a: douta_buf <= 22'h0000000000000000000000;
                12'h0e3b: douta_buf <= 22'h0000000000000000000000;
                12'h0e3c: douta_buf <= 22'h0000000000000000000000;
                12'h0e3d: douta_buf <= 22'h0000000000000000000000;
                12'h0e3e: douta_buf <= 22'h0000000000000000000000;
                12'h0e3f: douta_buf <= 22'h0000000000000000000000;
                12'h0e40: douta_buf <= 22'h0000000000000000000000;
                12'h0e41: douta_buf <= 22'h0000000000000000000000;
                12'h0e42: douta_buf <= 22'h0000000000000000000000;
                12'h0e43: douta_buf <= 22'h0000000000000000000000;
                12'h0e44: douta_buf <= 22'h0000000000000000000000;
                12'h0e45: douta_buf <= 22'h0000000000000000000000;
                12'h0e46: douta_buf <= 22'h0000000000000000000000;
                12'h0e47: douta_buf <= 22'h0000000000000000000000;
                12'h0e48: douta_buf <= 22'h0000000000000000000000;
                12'h0e49: douta_buf <= 22'h0000000000000000000000;
                12'h0e4a: douta_buf <= 22'h0000000000000000000000;
                12'h0e4b: douta_buf <= 22'h0000000000000000000000;
                12'h0e4c: douta_buf <= 22'h0000000000000000000000;
                12'h0e4d: douta_buf <= 22'h0000000000000000000000;
                12'h0e4e: douta_buf <= 22'h0000000000000000000000;
                12'h0e4f: douta_buf <= 22'h0000000000000000000000;
                12'h0e50: douta_buf <= 22'h0000000000000000000000;
                12'h0e51: douta_buf <= 22'h0000000000000000000000;
                12'h0e52: douta_buf <= 22'h0000000000000000000000;
                12'h0e53: douta_buf <= 22'h0000000000000000000000;
                12'h0e54: douta_buf <= 22'h0000000000000000000000;
                12'h0e55: douta_buf <= 22'h0000000000000000000000;
                12'h0e56: douta_buf <= 22'h0000000000000000000000;
                12'h0e57: douta_buf <= 22'h0000000000000000000000;
                12'h0e58: douta_buf <= 22'h0000000000000000000000;
                12'h0e59: douta_buf <= 22'h0000000000000000000000;
                12'h0e5a: douta_buf <= 22'h0000000000000000000000;
                12'h0e5b: douta_buf <= 22'h0000000000000000000000;
                12'h0e5c: douta_buf <= 22'h0000000000000000000000;
                12'h0e5d: douta_buf <= 22'h0000000000000000000000;
                12'h0e5e: douta_buf <= 22'h0000000000000000000000;
                12'h0e5f: douta_buf <= 22'h0000000000000000000000;
                12'h0e60: douta_buf <= 22'h0000000000000000000000;
                12'h0e61: douta_buf <= 22'h0000000000000000000000;
                12'h0e62: douta_buf <= 22'h0000000000000000000000;
                12'h0e63: douta_buf <= 22'h0000000000000000000000;
                12'h0e64: douta_buf <= 22'h0000000000000000000000;
                12'h0e65: douta_buf <= 22'h0000000000000000000000;
                12'h0e66: douta_buf <= 22'h0000000000000000000000;
                12'h0e67: douta_buf <= 22'h0000000000000000000000;
                12'h0e68: douta_buf <= 22'h0000000000000000000000;
                12'h0e69: douta_buf <= 22'h0000000000000000000000;
                12'h0e6a: douta_buf <= 22'h0000000000000000000000;
                12'h0e6b: douta_buf <= 22'h0000000000000000000000;
                12'h0e6c: douta_buf <= 22'h0000000000000000000000;
                12'h0e6d: douta_buf <= 22'h0000000000000000000000;
                12'h0e6e: douta_buf <= 22'h0000000000000000000000;
                12'h0e6f: douta_buf <= 22'h0000000000000000000000;
                12'h0e70: douta_buf <= 22'h0000000000000000000000;
                12'h0e71: douta_buf <= 22'h0000000000000000000000;
                12'h0e72: douta_buf <= 22'h0000000000000000000000;
                12'h0e73: douta_buf <= 22'h0000000000000000000000;
                12'h0e74: douta_buf <= 22'h0000000000000000000000;
                12'h0e75: douta_buf <= 22'h0000000000000000000000;
                12'h0e76: douta_buf <= 22'h0000000000000000000000;
                12'h0e77: douta_buf <= 22'h0000000000000000000000;
                12'h0e78: douta_buf <= 22'h0000000000000000000000;
                12'h0e79: douta_buf <= 22'h0000000000000000000000;
                12'h0e7a: douta_buf <= 22'h0000000000000000000000;
                12'h0e7b: douta_buf <= 22'h0000000000000000000000;
                12'h0e7c: douta_buf <= 22'h0000000000000000000000;
                12'h0e7d: douta_buf <= 22'h0000000000000000000000;
                12'h0e7e: douta_buf <= 22'h0000000000000000000000;
                12'h0e7f: douta_buf <= 22'h0000000000000000000000;
                12'h0e80: douta_buf <= 22'h0000000000000000000000;
                12'h0e81: douta_buf <= 22'h0000000000000000000000;
                12'h0e82: douta_buf <= 22'h0000000000000000000000;
                12'h0e83: douta_buf <= 22'h0000000000000000000000;
                12'h0e84: douta_buf <= 22'h0000000000000000000000;
                12'h0e85: douta_buf <= 22'h0000000000000000000000;
                12'h0e86: douta_buf <= 22'h0000000000000000000000;
                12'h0e87: douta_buf <= 22'h0000000000000000000000;
                12'h0e88: douta_buf <= 22'h0000000000000000000000;
                12'h0e89: douta_buf <= 22'h0000000000000000000000;
                12'h0e8a: douta_buf <= 22'h0000000000000000000000;
                12'h0e8b: douta_buf <= 22'h0000000000000000000000;
                12'h0e8c: douta_buf <= 22'h0000000000000000000000;
                12'h0e8d: douta_buf <= 22'h0000000000000000000000;
                12'h0e8e: douta_buf <= 22'h0000000000000000000000;
                12'h0e8f: douta_buf <= 22'h0000000000000000000000;
                12'h0e90: douta_buf <= 22'h0000000000000000000000;
                12'h0e91: douta_buf <= 22'h0000000000000000000000;
                12'h0e92: douta_buf <= 22'h0000000000000000000000;
                12'h0e93: douta_buf <= 22'h0000000000000000000000;
                12'h0e94: douta_buf <= 22'h0000000000000000000000;
                12'h0e95: douta_buf <= 22'h0000000000000000000000;
                12'h0e96: douta_buf <= 22'h0000000000000000000000;
                12'h0e97: douta_buf <= 22'h0000000000000000000000;
                12'h0e98: douta_buf <= 22'h0000000000000000000000;
                12'h0e99: douta_buf <= 22'h0000000000000000000000;
                12'h0e9a: douta_buf <= 22'h0000000000000000000000;
                12'h0e9b: douta_buf <= 22'h0000000000000000000000;
                12'h0e9c: douta_buf <= 22'h0000000000000000000000;
                12'h0e9d: douta_buf <= 22'h0000000000000000000000;
                12'h0e9e: douta_buf <= 22'h0000000000000000000000;
                12'h0e9f: douta_buf <= 22'h0000000000000000000000;
                12'h0ea0: douta_buf <= 22'h0000000000000000000000;
                12'h0ea1: douta_buf <= 22'h0000000000000000000000;
                12'h0ea2: douta_buf <= 22'h0000000000000000000000;
                12'h0ea3: douta_buf <= 22'h0000000000000000000000;
                12'h0ea4: douta_buf <= 22'h0000000000000000000000;
                12'h0ea5: douta_buf <= 22'h0000000000000000000000;
                12'h0ea6: douta_buf <= 22'h0000000000000000000000;
                12'h0ea7: douta_buf <= 22'h0000000000000000000000;
                12'h0ea8: douta_buf <= 22'h0000000000000000000000;
                12'h0ea9: douta_buf <= 22'h0000000000000000000000;
                12'h0eaa: douta_buf <= 22'h0000000000000000000000;
                12'h0eab: douta_buf <= 22'h0000000000000000000000;
                12'h0eac: douta_buf <= 22'h0000000000000000000000;
                12'h0ead: douta_buf <= 22'h0000000000000000000000;
                12'h0eae: douta_buf <= 22'h0000000000000000000000;
                12'h0eaf: douta_buf <= 22'h0000000000000000000000;
                12'h0eb0: douta_buf <= 22'h0000000000000000000000;
                12'h0eb1: douta_buf <= 22'h0000000000000000000000;
                12'h0eb2: douta_buf <= 22'h0000000000000000000000;
                12'h0eb3: douta_buf <= 22'h0000000000000000000000;
                12'h0eb4: douta_buf <= 22'h0000000000000000000000;
                12'h0eb5: douta_buf <= 22'h0000000000000000000000;
                12'h0eb6: douta_buf <= 22'h0000000000000000000000;
                12'h0eb7: douta_buf <= 22'h0000000000000000000000;
                12'h0eb8: douta_buf <= 22'h0000000000000000000000;
                12'h0eb9: douta_buf <= 22'h0000000000000000000000;
                12'h0eba: douta_buf <= 22'h0000000000000000000000;
                12'h0ebb: douta_buf <= 22'h0000000000000000000000;
                12'h0ebc: douta_buf <= 22'h0000000000000000000000;
                12'h0ebd: douta_buf <= 22'h0000000000000000000000;
                12'h0ebe: douta_buf <= 22'h0000000000000000000000;
                12'h0ebf: douta_buf <= 22'h0000000000000000000000;
                12'h0ec0: douta_buf <= 22'h0000000000000000000000;
                12'h0ec1: douta_buf <= 22'h0000000000000000000000;
                12'h0ec2: douta_buf <= 22'h0000000000000000000000;
                12'h0ec3: douta_buf <= 22'h0000000000000000000000;
                12'h0ec4: douta_buf <= 22'h0000000000000000000000;
                12'h0ec5: douta_buf <= 22'h0000000000000000000000;
                12'h0ec6: douta_buf <= 22'h0000000000000000000000;
                12'h0ec7: douta_buf <= 22'h0000000000000000000000;
                12'h0ec8: douta_buf <= 22'h0000000000000000000000;
                12'h0ec9: douta_buf <= 22'h0000000000000000000000;
                12'h0eca: douta_buf <= 22'h0000000000000000000000;
                12'h0ecb: douta_buf <= 22'h0000000000000000000000;
                12'h0ecc: douta_buf <= 22'h0000000000000000000000;
                12'h0ecd: douta_buf <= 22'h0000000000000000000000;
                12'h0ece: douta_buf <= 22'h0000000000000000000000;
                12'h0ecf: douta_buf <= 22'h0000000000000000000000;
                12'h0ed0: douta_buf <= 22'h0000000000000000000000;
                12'h0ed1: douta_buf <= 22'h0000000000000000000000;
                12'h0ed2: douta_buf <= 22'h0000000000000000000000;
                12'h0ed3: douta_buf <= 22'h0000000000000000000000;
                12'h0ed4: douta_buf <= 22'h0000000000000000000000;
                12'h0ed5: douta_buf <= 22'h0000000000000000000000;
                12'h0ed6: douta_buf <= 22'h0000000000000000000000;
                12'h0ed7: douta_buf <= 22'h0000000000000000000000;
                12'h0ed8: douta_buf <= 22'h0000000000000000000000;
                12'h0ed9: douta_buf <= 22'h0000000000000000000000;
                12'h0eda: douta_buf <= 22'h0000000000000000000000;
                12'h0edb: douta_buf <= 22'h0000000000000000000000;
                12'h0edc: douta_buf <= 22'h0000000000000000000000;
                12'h0edd: douta_buf <= 22'h0000000000000000000000;
                12'h0ede: douta_buf <= 22'h0000000000000000000000;
                12'h0edf: douta_buf <= 22'h0000000000000000000000;
                12'h0ee0: douta_buf <= 22'h0000000000000000000000;
                12'h0ee1: douta_buf <= 22'h0000000000000000000000;
                12'h0ee2: douta_buf <= 22'h0000000000000000000000;
                12'h0ee3: douta_buf <= 22'h0000000000000000000000;
                12'h0ee4: douta_buf <= 22'h0000000000000000000000;
                12'h0ee5: douta_buf <= 22'h0000000000000000000000;
                12'h0ee6: douta_buf <= 22'h0000000000000000000000;
                12'h0ee7: douta_buf <= 22'h0000000000000000000000;
                12'h0ee8: douta_buf <= 22'h0000000000000000000000;
                12'h0ee9: douta_buf <= 22'h0000000000000000000000;
                12'h0eea: douta_buf <= 22'h0000000000000000000000;
                12'h0eeb: douta_buf <= 22'h0000000000000000000000;
                12'h0eec: douta_buf <= 22'h0000000000000000000000;
                12'h0eed: douta_buf <= 22'h0000000000000000000000;
                12'h0eee: douta_buf <= 22'h0000000000000000000000;
                12'h0eef: douta_buf <= 22'h0000000000000000000000;
                12'h0ef0: douta_buf <= 22'h0000000000000000000000;
                12'h0ef1: douta_buf <= 22'h0000000000000000000000;
                12'h0ef2: douta_buf <= 22'h0000000000000000000000;
                12'h0ef3: douta_buf <= 22'h0000000000000000000000;
                12'h0ef4: douta_buf <= 22'h0000000000000000000000;
                12'h0ef5: douta_buf <= 22'h0000000000000000000000;
                12'h0ef6: douta_buf <= 22'h0000000000000000000000;
                12'h0ef7: douta_buf <= 22'h0000000000000000000000;
                12'h0ef8: douta_buf <= 22'h0000000000000000000000;
                12'h0ef9: douta_buf <= 22'h0000000000000000000000;
                12'h0efa: douta_buf <= 22'h0000000000000000000000;
                12'h0efb: douta_buf <= 22'h0000000000000000000000;
                12'h0efc: douta_buf <= 22'h0000000000000000000000;
                12'h0efd: douta_buf <= 22'h0000000000000000000000;
                12'h0efe: douta_buf <= 22'h0000000000000000000000;
                12'h0eff: douta_buf <= 22'h0000000000000000000000;
                12'h0f00: douta_buf <= 22'h0000000000000000000000;
                12'h0f01: douta_buf <= 22'h0000000000000000000000;
                12'h0f02: douta_buf <= 22'h0000000000000000000000;
                12'h0f03: douta_buf <= 22'h0000000000000000000000;
                12'h0f04: douta_buf <= 22'h0000000000000000000000;
                12'h0f05: douta_buf <= 22'h0000000000000000000000;
                12'h0f06: douta_buf <= 22'h0000000000000000000000;
                12'h0f07: douta_buf <= 22'h0000000000000000000000;
                12'h0f08: douta_buf <= 22'h0000000000000000000000;
                12'h0f09: douta_buf <= 22'h0000000000000000000000;
                12'h0f0a: douta_buf <= 22'h0000000000000000000000;
                12'h0f0b: douta_buf <= 22'h0000000000000000000000;
                12'h0f0c: douta_buf <= 22'h0000000000000000000000;
                12'h0f0d: douta_buf <= 22'h0000000000000000000000;
                12'h0f0e: douta_buf <= 22'h0000000000000000000000;
                12'h0f0f: douta_buf <= 22'h0000000000000000000000;
                12'h0f10: douta_buf <= 22'h0000000000000000000000;
                12'h0f11: douta_buf <= 22'h0000000000000000000000;
                12'h0f12: douta_buf <= 22'h0000000000000000000000;
                12'h0f13: douta_buf <= 22'h0000000000000000000000;
                12'h0f14: douta_buf <= 22'h0000000000000000000000;
                12'h0f15: douta_buf <= 22'h0000000000000000000000;
                12'h0f16: douta_buf <= 22'h0000000000000000000000;
                12'h0f17: douta_buf <= 22'h0000000000000000000000;
                12'h0f18: douta_buf <= 22'h0000000000000000000000;
                12'h0f19: douta_buf <= 22'h0000000000000000000000;
                12'h0f1a: douta_buf <= 22'h0000000000000000000000;
                12'h0f1b: douta_buf <= 22'h0000000000000000000000;
                12'h0f1c: douta_buf <= 22'h0000000000000000000000;
                12'h0f1d: douta_buf <= 22'h0000000000000000000000;
                12'h0f1e: douta_buf <= 22'h0000000000000000000000;
                12'h0f1f: douta_buf <= 22'h0000000000000000000000;
                12'h0f20: douta_buf <= 22'h0000000000000000000000;
                12'h0f21: douta_buf <= 22'h0000000000000000000000;
                12'h0f22: douta_buf <= 22'h0000000000000000000000;
                12'h0f23: douta_buf <= 22'h0000000000000000000000;
                12'h0f24: douta_buf <= 22'h0000000000000000000000;
                12'h0f25: douta_buf <= 22'h0000000000000000000000;
                12'h0f26: douta_buf <= 22'h0000000000000000000000;
                12'h0f27: douta_buf <= 22'h0000000000000000000000;
                12'h0f28: douta_buf <= 22'h0000000000000000000000;
                12'h0f29: douta_buf <= 22'h0000000000000000000000;
                12'h0f2a: douta_buf <= 22'h0000000000000000000000;
                12'h0f2b: douta_buf <= 22'h0000000000000000000000;
                12'h0f2c: douta_buf <= 22'h0000000000000000000000;
                12'h0f2d: douta_buf <= 22'h0000000000000000000000;
                12'h0f2e: douta_buf <= 22'h0000000000000000000000;
                12'h0f2f: douta_buf <= 22'h0000000000000000000000;
                12'h0f30: douta_buf <= 22'h0000000000000000000000;
                12'h0f31: douta_buf <= 22'h0000000000000000000000;
                12'h0f32: douta_buf <= 22'h0000000000000000000000;
                12'h0f33: douta_buf <= 22'h0000000000000000000000;
                12'h0f34: douta_buf <= 22'h0000000000000000000000;
                12'h0f35: douta_buf <= 22'h0000000000000000000000;
                12'h0f36: douta_buf <= 22'h0000000000000000000000;
                12'h0f37: douta_buf <= 22'h0000000000000000000000;
                12'h0f38: douta_buf <= 22'h0000000000000000000000;
                12'h0f39: douta_buf <= 22'h0000000000000000000000;
                12'h0f3a: douta_buf <= 22'h0000000000000000000000;
                12'h0f3b: douta_buf <= 22'h0000000000000000000000;
                12'h0f3c: douta_buf <= 22'h0000000000000000000000;
                12'h0f3d: douta_buf <= 22'h0000000000000000000000;
                12'h0f3e: douta_buf <= 22'h0000000000000000000000;
                12'h0f3f: douta_buf <= 22'h0000000000000000000000;
                12'h0f40: douta_buf <= 22'h0000000000000000000000;
                12'h0f41: douta_buf <= 22'h0000000000000000000000;
                12'h0f42: douta_buf <= 22'h0000000000000000000000;
                12'h0f43: douta_buf <= 22'h0000000000000000000000;
                12'h0f44: douta_buf <= 22'h0000000000000000000000;
                12'h0f45: douta_buf <= 22'h0000000000000000000000;
                12'h0f46: douta_buf <= 22'h0000000000000000000000;
                12'h0f47: douta_buf <= 22'h0000000000000000000000;
                12'h0f48: douta_buf <= 22'h0000000000000000000000;
                12'h0f49: douta_buf <= 22'h0000000000000000000000;
                12'h0f4a: douta_buf <= 22'h0000000000000000000000;
                12'h0f4b: douta_buf <= 22'h0000000000000000000000;
                12'h0f4c: douta_buf <= 22'h0000000000000000000000;
                12'h0f4d: douta_buf <= 22'h0000000000000000000000;
                12'h0f4e: douta_buf <= 22'h0000000000000000000000;
                12'h0f4f: douta_buf <= 22'h0000000000000000000000;
                12'h0f50: douta_buf <= 22'h0000000000000000000000;
                12'h0f51: douta_buf <= 22'h0000000000000000000000;
                12'h0f52: douta_buf <= 22'h0000000000000000000000;
                12'h0f53: douta_buf <= 22'h0000000000000000000000;
                12'h0f54: douta_buf <= 22'h0000000000000000000000;
                12'h0f55: douta_buf <= 22'h0000000000000000000000;
                12'h0f56: douta_buf <= 22'h0000000000000000000000;
                12'h0f57: douta_buf <= 22'h0000000000000000000000;
                12'h0f58: douta_buf <= 22'h0000000000000000000000;
                12'h0f59: douta_buf <= 22'h0000000000000000000000;
                12'h0f5a: douta_buf <= 22'h0000000000000000000000;
                12'h0f5b: douta_buf <= 22'h0000000000000000000000;
                12'h0f5c: douta_buf <= 22'h0000000000000000000000;
                12'h0f5d: douta_buf <= 22'h0000000000000000000000;
                12'h0f5e: douta_buf <= 22'h0000000000000000000000;
                12'h0f5f: douta_buf <= 22'h0000000000000000000000;
                12'h0f60: douta_buf <= 22'h0000000000000000000000;
                12'h0f61: douta_buf <= 22'h0000000000000000000000;
                12'h0f62: douta_buf <= 22'h0000000000000000000000;
                12'h0f63: douta_buf <= 22'h0000000000000000000000;
                12'h0f64: douta_buf <= 22'h0000000000000000000000;
                12'h0f65: douta_buf <= 22'h0000000000000000000000;
                12'h0f66: douta_buf <= 22'h0000000000000000000000;
                12'h0f67: douta_buf <= 22'h0000000000000000000000;
                12'h0f68: douta_buf <= 22'h0000000000000000000000;
                12'h0f69: douta_buf <= 22'h0000000000000000000000;
                12'h0f6a: douta_buf <= 22'h0000000000000000000000;
                12'h0f6b: douta_buf <= 22'h0000000000000000000000;
                12'h0f6c: douta_buf <= 22'h0000000000000000000000;
                12'h0f6d: douta_buf <= 22'h0000000000000000000000;
                12'h0f6e: douta_buf <= 22'h0000000000000000000000;
                12'h0f6f: douta_buf <= 22'h0000000000000000000000;
                12'h0f70: douta_buf <= 22'h0000000000000000000000;
                12'h0f71: douta_buf <= 22'h0000000000000000000000;
                12'h0f72: douta_buf <= 22'h0000000000000000000000;
                12'h0f73: douta_buf <= 22'h0000000000000000000000;
                12'h0f74: douta_buf <= 22'h0000000000000000000000;
                12'h0f75: douta_buf <= 22'h0000000000000000000000;
                12'h0f76: douta_buf <= 22'h0000000000000000000000;
                12'h0f77: douta_buf <= 22'h0000000000000000000000;
                12'h0f78: douta_buf <= 22'h0000000000000000000000;
                12'h0f79: douta_buf <= 22'h0000000000000000000000;
                12'h0f7a: douta_buf <= 22'h0000000000000000000000;
                12'h0f7b: douta_buf <= 22'h0000000000000000000000;
                12'h0f7c: douta_buf <= 22'h0000000000000000000000;
                12'h0f7d: douta_buf <= 22'h0000000000000000000000;
                12'h0f7e: douta_buf <= 22'h0000000000000000000000;
                12'h0f7f: douta_buf <= 22'h0000000000000000000000;
                12'h0f80: douta_buf <= 22'h0000000000000000000000;
                12'h0f81: douta_buf <= 22'h0000000000000000000000;
                12'h0f82: douta_buf <= 22'h0000000000000000000000;
                12'h0f83: douta_buf <= 22'h0000000000000000000000;
                12'h0f84: douta_buf <= 22'h0000000000000000000000;
                12'h0f85: douta_buf <= 22'h0000000000000000000000;
                12'h0f86: douta_buf <= 22'h0000000000000000000000;
                12'h0f87: douta_buf <= 22'h0000000000000000000000;
                12'h0f88: douta_buf <= 22'h0000000000000000000000;
                12'h0f89: douta_buf <= 22'h0000000000000000000000;
                12'h0f8a: douta_buf <= 22'h0000000000000000000000;
                12'h0f8b: douta_buf <= 22'h0000000000000000000000;
                12'h0f8c: douta_buf <= 22'h0000000000000000000000;
                12'h0f8d: douta_buf <= 22'h0000000000000000000000;
                12'h0f8e: douta_buf <= 22'h0000000000000000000000;
                12'h0f8f: douta_buf <= 22'h0000000000000000000000;
                12'h0f90: douta_buf <= 22'h0000000000000000000000;
                12'h0f91: douta_buf <= 22'h0000000000000000000000;
                12'h0f92: douta_buf <= 22'h0000000000000000000000;
                12'h0f93: douta_buf <= 22'h0000000000000000000000;
                12'h0f94: douta_buf <= 22'h0000000000000000000000;
                12'h0f95: douta_buf <= 22'h0000000000000000000000;
                12'h0f96: douta_buf <= 22'h0000000000000000000000;
                12'h0f97: douta_buf <= 22'h0000000000000000000000;
                12'h0f98: douta_buf <= 22'h0000000000000000000000;
                12'h0f99: douta_buf <= 22'h0000000000000000000000;
                12'h0f9a: douta_buf <= 22'h0000000000000000000000;
                12'h0f9b: douta_buf <= 22'h0000000000000000000000;
                12'h0f9c: douta_buf <= 22'h0000000000000000000000;
                12'h0f9d: douta_buf <= 22'h0000000000000000000000;
                12'h0f9e: douta_buf <= 22'h0000000000000000000000;
                12'h0f9f: douta_buf <= 22'h0000000000000000000000;
                12'h0fa0: douta_buf <= 22'h0000000000000000000000;
                12'h0fa1: douta_buf <= 22'h0000000000000000000000;
                12'h0fa2: douta_buf <= 22'h0000000000000000000000;
                12'h0fa3: douta_buf <= 22'h0000000000000000000000;
                12'h0fa4: douta_buf <= 22'h0000000000000000000000;
                12'h0fa5: douta_buf <= 22'h0000000000000000000000;
                12'h0fa6: douta_buf <= 22'h0000000000000000000000;
                12'h0fa7: douta_buf <= 22'h0000000000000000000000;
                12'h0fa8: douta_buf <= 22'h0000000000000000000000;
                12'h0fa9: douta_buf <= 22'h0000000000000000000000;
                12'h0faa: douta_buf <= 22'h0000000000000000000000;
                12'h0fab: douta_buf <= 22'h0000000000000000000000;
                12'h0fac: douta_buf <= 22'h0000000000000000000000;
                12'h0fad: douta_buf <= 22'h0000000000000000000000;
                12'h0fae: douta_buf <= 22'h0000000000000000000000;
                12'h0faf: douta_buf <= 22'h0000000000000000000000;
                12'h0fb0: douta_buf <= 22'h0000000000000000000000;
                12'h0fb1: douta_buf <= 22'h0000000000000000000000;
                12'h0fb2: douta_buf <= 22'h0000000000000000000000;
                12'h0fb3: douta_buf <= 22'h0000000000000000000000;
                12'h0fb4: douta_buf <= 22'h0000000000000000000000;
                12'h0fb5: douta_buf <= 22'h0000000000000000000000;
                12'h0fb6: douta_buf <= 22'h0000000000000000000000;
                12'h0fb7: douta_buf <= 22'h0000000000000000000000;
                12'h0fb8: douta_buf <= 22'h0000000000000000000000;
                12'h0fb9: douta_buf <= 22'h0000000000000000000000;
                12'h0fba: douta_buf <= 22'h0000000000000000000000;
                12'h0fbb: douta_buf <= 22'h0000000000000000000000;
                12'h0fbc: douta_buf <= 22'h0000000000000000000000;
                12'h0fbd: douta_buf <= 22'h0000000000000000000000;
                12'h0fbe: douta_buf <= 22'h0000000000000000000000;
                12'h0fbf: douta_buf <= 22'h0000000000000000000000;
                12'h0fc0: douta_buf <= 22'h0000000000000000000000;
                12'h0fc1: douta_buf <= 22'h0000000000000000000000;
                12'h0fc2: douta_buf <= 22'h0000000000000000000000;
                12'h0fc3: douta_buf <= 22'h0000000000000000000000;
                12'h0fc4: douta_buf <= 22'h0000000000000000000000;
                12'h0fc5: douta_buf <= 22'h0000000000000000000000;
                12'h0fc6: douta_buf <= 22'h0000000000000000000000;
                12'h0fc7: douta_buf <= 22'h0000000000000000000000;
                12'h0fc8: douta_buf <= 22'h0000000000000000000000;
                12'h0fc9: douta_buf <= 22'h0000000000000000000000;
                12'h0fca: douta_buf <= 22'h0000000000000000000000;
                12'h0fcb: douta_buf <= 22'h0000000000000000000000;
                12'h0fcc: douta_buf <= 22'h0000000000000000000000;
                12'h0fcd: douta_buf <= 22'h0000000000000000000000;
                12'h0fce: douta_buf <= 22'h0000000000000000000000;
                12'h0fcf: douta_buf <= 22'h0000000000000000000000;
                12'h0fd0: douta_buf <= 22'h0000000000000000000000;
                12'h0fd1: douta_buf <= 22'h0000000000000000000000;
                12'h0fd2: douta_buf <= 22'h0000000000000000000000;
                12'h0fd3: douta_buf <= 22'h0000000000000000000000;
                12'h0fd4: douta_buf <= 22'h0000000000000000000000;
                12'h0fd5: douta_buf <= 22'h0000000000000000000000;
                12'h0fd6: douta_buf <= 22'h0000000000000000000000;
                12'h0fd7: douta_buf <= 22'h0000000000000000000000;
                12'h0fd8: douta_buf <= 22'h0000000000000000000000;
                12'h0fd9: douta_buf <= 22'h0000000000000000000000;
                12'h0fda: douta_buf <= 22'h0000000000000000000000;
                12'h0fdb: douta_buf <= 22'h0000000000000000000000;
                12'h0fdc: douta_buf <= 22'h0000000000000000000000;
                12'h0fdd: douta_buf <= 22'h0000000000000000000000;
                12'h0fde: douta_buf <= 22'h0000000000000000000000;
                12'h0fdf: douta_buf <= 22'h0000000000000000000000;
                12'h0fe0: douta_buf <= 22'h0000000000000000000000;
                12'h0fe1: douta_buf <= 22'h0000000000000000000000;
                12'h0fe2: douta_buf <= 22'h0000000000000000000000;
                12'h0fe3: douta_buf <= 22'h0000000000000000000000;
                12'h0fe4: douta_buf <= 22'h0000000000000000000000;
                12'h0fe5: douta_buf <= 22'h0000000000000000000000;
                12'h0fe6: douta_buf <= 22'h0000000000000000000000;
                12'h0fe7: douta_buf <= 22'h0000000000000000000000;
                12'h0fe8: douta_buf <= 22'h0000000000000000000000;
                12'h0fe9: douta_buf <= 22'h0000000000000000000000;
                12'h0fea: douta_buf <= 22'h0000000000000000000000;
                12'h0feb: douta_buf <= 22'h0000000000000000000000;
                12'h0fec: douta_buf <= 22'h0000000000000000000000;
                12'h0fed: douta_buf <= 22'h0000000000000000000000;
                12'h0fee: douta_buf <= 22'h0000000000000000000000;
                12'h0fef: douta_buf <= 22'h0000000000000000000000;
                12'h0ff0: douta_buf <= 22'h0000000000000000000000;
                12'h0ff1: douta_buf <= 22'h0000000000000000000000;
                12'h0ff2: douta_buf <= 22'h0000000000000000000000;
                12'h0ff3: douta_buf <= 22'h0000000000000000000000;
                12'h0ff4: douta_buf <= 22'h0000000000000000000000;
                12'h0ff5: douta_buf <= 22'h0000000000000000000000;
                12'h0ff6: douta_buf <= 22'h0000000000000000000000;
                12'h0ff7: douta_buf <= 22'h0000000000000000000000;
                12'h0ff8: douta_buf <= 22'h0000000000000000000000;
                12'h0ff9: douta_buf <= 22'h0000000000000000000000;
                12'h0ffa: douta_buf <= 22'h0000000000000000000000;
                12'h0ffb: douta_buf <= 22'h0000000000000000000000;
                12'h0ffc: douta_buf <= 22'h0000000000000000000000;
                12'h0ffd: douta_buf <= 22'h0000000000000000000000;
                12'h0ffe: douta_buf <= 22'h0000000000000000000000;
                12'h0fff: douta_buf <= 22'h0000000000000000000000;
            endcase
        end
    end

    assign douta = douta_buf;
endmodule
